//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   2023 ICLAB Fall Course
//   Lab03      : BRIDGE
//   Author     : Ting-Yu Chang
//                
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : BRIDGE_encrypted.v
//   Module Name : BRIDGE
//   Release version : v1.0 (Release Date: Sep-2023)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

module BRIDGE(
    // Input Signals
    clk,
    rst_n,
    in_valid,
    direction,
    addr_dram,
    addr_sd,
    // Output Signals
    out_valid,
    out_data,
    // DRAM Signals
    AR_VALID, AR_ADDR, R_READY, AW_VALID, AW_ADDR, W_VALID, W_DATA, B_READY,
	AR_READY, R_VALID, R_RESP, R_DATA, AW_READY, W_READY, B_VALID, B_RESP,
    // SD Signals
    MISO,
    MOSI
);


`protected
HT&[\)&JSab@E5b;a\DRCd,K_RC&AEeeEJYOd1WNTF,(Z@\H(=M2.)IC4&<#>S8c
35ga&Q3JWeRBf_O[EM8;[A^F)f&>DbM#:$
`endprotected
input clk, rst_n;
input in_valid;
input direction;
input [12:0] addr_dram;
input [15:0] addr_sd;


`protected
K2:_W\NLaC+,fZ)[W?Fa]BJU+DagUdNI>@P\L7;-X2f?edY9egOL&)U6WO,TKHG6
9d@XGOHITH)?a@V(=?L:-<e4)OgebH9C;$
`endprotected
output reg out_valid;
output reg [7:0] out_data;


`protected
Za?^Bb0>)J;<.IFNSLO.YK/]H##X)-UE.:<I^e\gY4SI]S,FH<.W2)@B)ae&CfG0
;Q02GU<U)T?XdC^G7TOQ)?b4\GRF/<R3K<.\:VP[K.d4\7[ZaI6gZc^:?(D93UNeS$
`endprotected
output reg [31:0] AW_ADDR;
output reg AW_VALID;
input AW_READY;

`protected
b=ITgE;f)I2g7IQZ;H^Z9@/g].-^T,>7SF62AG4QLNH-Ka6Te,_O/)+V#+JL,^bR
<N3=]I0B_90(F^YAOKM&>=H;2)28efbS?$
`endprotected
output reg W_VALID;
output reg [63:0] W_DATA;
input W_READY;

`protected
5V09\W+]3;#:W+(E_SOEQR5gD+GIc/WK6]Z-9@Pg2&bD[AG)OI/D,))N8JU4Ng>A
aJ9V=TQ;/1-T8HV[3b+_La]AG_)L29LG,/&3N>O2F(TDC$
`endprotected
input B_VALID;
input [1:0] B_RESP;
output reg B_READY;

`protected
<DZT2_PL\&]Bg.S)<-UE6,CK1/6IZS;J59\6RC[K0]Q-QZ/X&HMW4)=A&TB.;1FH
CW3TZT57OL=A<((0E(]A-W;Q,[(>7cL91H#e(Nc=,a:-A$
`endprotected
output reg [31:0] AR_ADDR;
output reg AR_VALID;
input AR_READY;

`protected
eG2BD17VKJ/]HbbQdEVBQ@BP5ZT_eG?5;#,NFe3+?Fc?f@C7<0-W2)Q7AR/e0+G?
A_BP7^XLL1(A2MaH7R_)K)2Wd+4YTHY1>$
`endprotected
input [63:0] R_DATA;
input R_VALID;
input [1:0] R_RESP;
output reg R_READY;


`protected
0b=e\76gWF<D2<MP1?&GWe6GC\C6g0E_G?/ed;2D9R+]6M:4F)74-)>O]3TQHQR#
cQ+d5OGd8QN4\,)<=U4.7<6G7$
`endprotected
input MISO;
output reg MOSI;


`protected
(3dSZN;\G/U]:38gEO#\\:N1;UT34W7I(>B5de+^M\.c3-?HO_^X2)b+9RId]E[I
3AQI\Je=)\CW@>D35N<?g/5\@9WPI)Z\]c8gaN-^>@BA.f)N9F:I3CG6fYLI4^->
XFgMB5T:W9WXN53cT5DY.3V\;YXH.?I6MZ-[X80Ze6U49E7IAC:>^2gc&deQ)C96
1A[:3M<7+3-g\+=0F7B^bY5(O^f[>Ag#L&=2Z2,;-.S.S.GB021.P7^be:#7cJ&/
<.9e_2gE//]V/RY^S&fNcCD_g/0&;K.c198a?1de#&;[;(+C]C+#e_<MZYUU#9C>
dQLK]YNF=YU:88TLV7>c@_2,EJcOAg<,#eOb8cUW+8;)\3;38?b\J+Pf&HK3T+/-
I[&gTTXfI>?^S^fNT<AV@dG[2X>T9MYU>2b7Z2FID#K<JW[KU^=g[Y:YWC.C&S8U
;\D\X/C8WQJE-U\GgdT):2e]:K+5<D;?[Y+:SOdT4BbT_B=-ARL=&_L+TQcOC)1Y
//GgEb[e/T156cc\Le?@1Yc^&0]8AA(db8[:8O?J04>PTO+98S6D#B7PJRb@/>/T
+^_3N0\8<.A+66<7IK8C[46Y]/eP5Bf>G?3<3U3VBe0;Y=^JX[D)g.d2W?H_[c-^
3#.,aC1;ZUP9>^UZ,g)0[E\0Pf?+]=IW\f(g#;;4Q)9^R-I)ULOHZ0dGa>J)SWYg
FcC(UMJgDXd27Rg48cf>H(4N6D1]bM=QVe;<O#;ZO;W;3d)aLI+e<^>03[0[&8+3
S_7#MW6SW]aMBCeWIRB8Td>3^KcI?Kc@(PC_B7^^43f2OPLG+6+PeO:@>[6RJE+K
8M8g8#FRNO/+RPfdP<cTgbXA>eTY[&K&ac24P-92feO7:bdS@2O&X9]#K:ADb2Lg
Qbc4Zg-WJ-&19<XG\.A5]62PTSI0>5(-,Y-fVM>2-EgSeP7Pg-=WEd:JQ13?1M@0
.+4_WHaJ.G_(>g#-L#=/U[XcaL_G#PM-@9G>25&ZORI.4&E?G@([)T&0:e=aWA3E
GF9U9HDFb>)2G@A>9EJKY@-0aK(@RH=Pa5+_86a+(JDLQ(\00^H)[1Z4NcN,R:e1
P[LbLXBd#Hf+1EN4SaC@](_\QR9)gV;#X8Pe?7&H;+d5-><=HfMV\N8g\^&6#?FY
4\Ib9.gB#;S/E@R44PJ2D74ISO=94DF#WW(;RCM0F[WUI16cP^d_(9Ef0S#L\E6L
OCPSBOG1(S;E6J8E@RaVT;eKSf_E>QK5;_VRUJ5KbcLW+?6L9@Nd9-8aLL#f(8f6
:VJOE?B2IF^^0-4gE+7P>b#a+GNMZA?=]P>;S]E)FPQ>a\g#b/IJUA@L#NNfU#A>
@PAfW)IgZgYK(YIdd9:XFQYe8VA&PW>&.g>\@-g_Q>X>N>3=J._6EQVeg1\TD0ec
F/E[2U8)gXdW@_T;e)UFE1HA^2/T=ZHC6g(5;7e?_2+8NMWNZYE[A5VQ<d.UUF(_
6N5+_?abUH/6=3^_1(EAL<2P;5^KE&4M=JB@XR6(RXPfOUL3V]@)_Kd1.6,]G.c6
2>c+a/(_8\3GEWX>2&A=E]9->aU>dA(O6PKQ?ET(\-ZJbS=,gWc)]J(6CEYZ\#2B
[gL-AP3?ZBTEUHMeeg4>VZ9^B(bPXVCcD=3U<Rf2/#XXA6RZA&<DU&4FZ-]ZX6=f
N13dZ8^]@RB+NSPH1JedUA=9KZ\X](S)F_[>00]++[(\PE(BAY,<[C:d)3eSGe:5
H^N+g;#U4/7<0K<\X_MfWC(1Vg0V2-dGYIDb.YXC64dNFN6+VDD)@T5E[5RL;dT[
=:2E2YcVM/(ab05Y2T=?5YTeEHCKSM^5K55N;cC.;R08N,BU1U]T,UI08-Cf_SFE
7aR:aJg[H8DQQ.[Y)9)/+d+ZIc)N>P6g.6TO&6U_aG+B\Xb1<P?YDD3K9J>M)Ffe
R_+E-S-MFf6I,I./cZHb]Tb2IEWg+-:M@@1PEFNdKF[_QP9I<&E_NP43ac1;EW^)
_YLN18f8HCcWeNL/,\9E=TSULZD(.WUZ-,F>C)G@F).A/Ge+WL8aNCTRg10KHEaL
<[BfO@2KLP2b9c+g55fM26afe9Yg6R=B\E(&<22N@=0C,,MB8IeR7@Pe\PG:++JW
6#Dc7AVX#(O?.&YPJf^=81X[C8@ZQ_ZX-O[Q8NTcdd:HX)N]d<UcUP#T>,J4.BT7
_eSC@^SX2JH,&dGaL0c27T]R@Ce11M>^.1f7JI761MUJ[d_Mf>N&+[2<\G&U^AeU
\YQ/YKEH.;ICJ.:-NbHG^E.T(.:[U1K__+1UZVEg+^30#X/,L3ag_]+.4C4Y?@Z[
CHGNK8,V7<e5cgJ-9X6I>V-.7NW(+4;6G,+&[=@/,:8WR#a_XWRH-A&:0&?bRMb6
B^UI];/[g@@?(#\OaYI0YgNJT[ZR6cE/V1N6<8g9#UO7AD&VMg4WJVe(IF\IBgAF
3Y.9L8a,O0>7?:,+,M8OC,]INDQ>7VY3S^\aVbK13SQ)5g;RZJ.^9B92>TSI&f_4
5OAX@fQeWLL]\9C>,\2/+edaZ,NG3c5QaDINE[<.L69H:6).H1#?S5JNWe4DKB,V
_<Pg5&_]]B@<FZRd<.=_g64?T0=_[KGC6g<L=BHSOH&L6\Jf;6+Jg.F/2,UeV,.T
&;\UdX/_>6OK5S6PIfA1,IR(WEC:Z(MDa^N]]\HK=]A<gfCDbWd_aX44&J/G&WKT
b+ZPfc:S&Q7_:NI1=2N81C>F4OD-Xa<#W1YV<\3<AVUdBWS?G+_;BZP[>LgaMF4+
5[Q=.^:,QFM6-)a@I.UPD;A+S:M.0Y#IZ^f,9ME,;P5>3F>gVJe#DFNcEH#IQ\DY
-ZD_JG,QB.D]fOA1dUUISF+X[g?P+1A,Ye\1E(7#?Kg,_PJ9bR??MA[I)^=#-ONM
/PVR-95NBIPM2G@c,+:SBS1R#fF0KH#:a09M8/D)H/HcfVEE;.ME[^>OK#/KI:3M
;LFCR9-O&M+T0bGB@WULGO\2e/8#Q#D,_N#?d5_PDX2d-8GYSW3a2J>)IMUX;:JW
KdRf<UD>+UEZBZcfga3F)fL?[57?=E^LT@c_\:P]dO5@/1cNT,Y,BgANK=-CR/Of
AUIZgVfEf4>->T^2ERgeGc,cBSPRS1_J;L6a8_8L:HJ_/WX(BdWERRJ6211U4[:?
FQf-@89F+1@63XU[^6E;H^ZU6?W<5X?YZX28>]Q)=U:ATV+(Y,\J5VBK^Q/#g741
Ec8&AJGYX]9R_PS-Z_1#,U02.Y#W^&-eT0^.^G+dJ(A_7(R,CT>&HN-^L#f1bHOb
aK0^&4\/AOc7C)S^NPD7VRXXcGbC2Z/?-V[3+K+R]P/7KPd+?:9I&@5OaD_d8M6?
C]9;SS6#ZV[c&1]98:d.Q,g)D^DQC3E\MK]>\ODRAS6L+dH(-H[XB9=(AJMAPSK]
&1B:6gI++FIT+OPZeV(J\Cb=W2#6^R286W8CL3X0OO=CU^a.EO=Og2+b62HQ,PdQ
XC/+70F//J^58\^4PYgJO8A8^cJUFGgG@V)]7gW3]#XN\ZN\(2K.M_1G=9TaS9NX
Tb&N:+g7NGOG-C#_#=X8(^4OV9O39TM9@K(LddZdgWD5Fc)I//CMD1Q4I->?g/R?
\c5K/946SMG5K&Q=OAb]RP7P+d^>W7gJACb#3=IP170^J/:Q2SgF;#Yc2E0EN?(L
+Pe1DV&?K5Z;224f_@AX\@E67IgPda6L0b;#bL(c.Fab5GS?8V_&De)>/f6f]11)
4>;A^[LegB0_:];(TKJ/Z5OVU,@cQ\VU\e1bPe98N.^:8\9ON,]b]R-.bR]N^5C3
RYg(11KVA6WJV]\86LC9->XM>baI=U<(d12f;>CB[1--2c<0Pb>IAb,&bFW;KfD(
PFf-XB87<[FP9RNgK,^)G@J6=bPKW:;CCAPV<bV.K&b:EM/W/6MVH]MaW<2#?BN_
[2#-PcSKX70]D@-=:Z>+0aZ6LQ,gd-8YYO#fO)S>)1Q-@c?5U@c7b9/AHNIA[QPK
P8/3:)DA-R/d6A/.];a\Xb;6>a?#>?dNK5U\fOe-S?M^Z5^,F\/9cWP,.?gVP[4L
g2])S\gG&AP.@YbV]bH<H\g-857X,S8SR;JEJ9G0[@B@2WKT>YgNC[(fZfcF=3-Y
SbM=W/O4>Ae.SfXBVg8)=L:bN?Wa,/,b+2+^:VgedLa9/FQYOV-JR3O:D^0YCIIU
?b+OgU)QE&_&__RZA0V&>Cb64<Z5-M7PZfPZ;TQ0(S5-CH\L;WC<Qg8U#GY;TVPI
9.JLGdLc#VdBU,gbH-827)=&O5KD=b4:5NXd0+7\>1]A?U&1(S5II5E&&A-1d/[6
eRBNW1A]_f<.&feSJLX-a&5P8+TXa9A1L1>1=93/LG/[bWUT?bb1L09KCEa0V\]Z
:aR8)Jd(C?4#/4;U<G(7FI4K)O3R^:J0]@=H^M[+6b)@UEVbRSIHUNWYNfSXQ@-9
NeWLe)+;+A@77]BN)D5a#BF6=:YcHfX=<S[BDJ\Zd+A8H0-1UH8:XE.:a97(5RbE
I\[RLTGWCA4_,AQ^2EKfC-3/AXJB6Y)O<^57-37<D=NX/931b-.Y8>8c(5BMQ;J:
+Y&?e&D817A@S.?A(>=AOB3KD/;L=&E>])>Q59H_a?bRYMMY.XHMDZFb4.5UT/.N
,bTJ?5+Q;9,LHY2FBV&YY3X:6B=-6d@W+337&&(50cN)<O8,Fa<S.TeLQC6<Y5fL
Y4:I&N1Z535EYIIeZ?HeO0G:eW,THb)JY2A_Sb1gRRT._\&Q<[1[)</b^<AHT@ff
]#?XR^1cJ#E9YS5,7(UeYI^d/UIB7?L[Qd(5:JJe6/P9;PH+^Q=@-^CE9dZ,GB^e
WFC1]5Y6Z#-f33d\+,39V6/,Y\BVMg_75,R3=6J[Ne;FO;G.HXV9QM8\X]#;+ed7
IM&MbEB7-87\DM(91C/6AVM>G(aPbAEM<T5-=G9I^RON7D<LHE/48cgA+V]fc?R,
.([H@cIGZSI2CH3?\2YZ5Xc_Oc8.RO#=f=@;0G/;fQ4T_BAf+@VG5Z0V)WOX#K78
^b-gVd;&,KNVU9AIC<g>f85A\5Yd5d(fB#8NHY#FX4+2a;O(EFc=#(FDJbJg_\^a
Q5>^YcWN9(DAA[I)._RD[3WcA8N.Qc[.2([SP59WL?]@K)3ICgBL<a;(3O4#4PfF
B?U\@F(d:&AV>VAO[QA=f1P:ZdB+/dC]d:1H14DTb9HW+@S(c5M.(]C+]LYRG640
gF/B#L1Q&U2Q<;9c34^35G6TKffNMa5HW4I49&FC57W-7T9J9J1^^<^Yd5X&OQeX
e]:D)HJH9Z7A(9R;?YDaI9EK6<#<81_=]J&JB;,7@QU5Uc+LEQTVD6,fCO<c]H+D
JOFQJX-BA?6QV35GWM=<FNgQE+WT1gV:c)5/@3<H:P74g1/Q[c0=EZ7H@cX7B+S8
-DF;)<].]Ud&a)fU.^f9_.,d/WbR1KPfT_9KO.19eI@MG[?b+3b?QAYb,.06ddbd
b#?PNSN]PJbT-fCI2EZ_YM/27fZU5OJKS5=b4I42AbGbZVOFD@7AT,A0<UgG1GGS
2Pc?JH/;^#UA)O[B[.Ud/OE(>5(11G.1N>0TA,RRMZe=9BdLW/WU#gIQ/f42.1X1
P<PG(Bb>8]<NE<>JZ[KWCAFI,.02.7Q.^1g5V-GNE:DR33#4aBOPb2IK9TJ71E;,
KL@?=\[SS:(R-=&]1WB(Cc.-6ECF.ZV@UG>P)[7PH0[e1KW_6^^O:Q9D4L4F?CdK
KBIEEMaXJ#Ma_Aa6:N2RICZ^#7@HF],fI,BfX7RG?XAbUe<^:E04YL@)YV5-<B.B
KGCKQg[BPR6Dgf:BK]))A]If:B]fO&@c(AB]G=UD&5g5[L[=YT+aUS?,K)b-TQ)W
^?0]&\;^[g5>L.JLIO5bK1A(<AHI77b7K?_fgYOa3&W..Ug=UJ_aQ,)HV_9O]0#C
U6MD7<WT5R>P?FCU>;V1K6)R>+6:Jd9V=.^,^QQ+AY?CQcU8BRVUN1?3.)K#WfZQ
L^Vb>3LYVKOORH-f=1\FUPZP3Ld-a.EQI6NgM5\S):YQ=D,J6H&Cf8aS#;g,)ae7
3UP72W6EE4==a^5KeQ6\cgBPW^G?89-8e6SYU@^@@J88IA4aLJc.:=Ef+f^;C;&d
-<^W@V=R6ZC5/_8IJMW3KaNXV,^2YA&QN[>_,K)J7US=DHg@1P.V3>&;DfF=Ma&[
Z7S<R,d?803A[c3@J__M@2]W3E4Ag7;>>0TUDfPa4Z(=_9MSeNA>KSW/LPN[MI^Y
.P#PG?DI:D@[d,_P,L47\=(86:?.SV2@PQ_Z#+NbSXTZ:-&QV\dINg.6;.Pef/HT
:8B(g6T+:EgcTKKUd&[CNID#])D<#2Vg0/TRXZKdA=51T=&IERAbc#T:MISf8O9]
?dYIIegc@Nc2=dcKXDYQ)gI_aa_MFWDg52R8#ZQ>[7&+^DZgFdg+[?SBTLgTV)?(
S[PCRD9d_DcVHb_#/>Y7>U)&3,Ld974R=:bV&GPSCe[OBeO1>&S)K2</?VGQ&Df#
Ma0>VADd<VBK:CL1#^Q+,#[aLe,>VY\J8MNKa=FISfE\K;eU#HV?Y8/[2/)]ge?Y
=DQP6Z=aL-EPfKRa[&gD1ZS3;(V8Sd5>1/<+R@:L87<Yb86N3,J[Q7d&g1c,N3fG
\0Tf]MbD8<6&I9(a28c]C9>S5eN8Q53]I90T#4_bME5J7@ATbZ3Fd].SQ)ZY[=)<
8RGaR(cH4+)a1EA-?D2/W(7ZB-babbF>Ea5FaOEgDC#Yc46]0LRX)c&.;2Y=KX\#
;\C][B;LSHQ)f,L7@7bLcT8/L\Rfcd(OJf/2YQ-7CB,U)VW5&e9O>C^\_MebR4[E
c;Db_e?ECD[P,3K[@WG@N]>)(C6TZ,g<[@ALSVOJI=</UReA=#/18Z]5K8/K76_X
E,5QE<[Q\.@SH+2cX))UQMQHS,6[H/+:fg:CNJ[FLPfC3T7AeAY@TSF_&&@3A5TI
@W&I=;F.A#6.J5R\H/RR05MM+[=^XaF;F(H&gJ\G-c70LZIdP1O6S?6PVEKK@>Y4
OCUaGK,UGf#(60X;.N&)8XY<eb/3T52-AIcCTdVG,aN\RYec_W\)[(D#e/c5WV6A
[2ALf#&7#dcb.6\;[U6H<[1#@\,^<a0M(&e@U,\P?XZR>_9SZ(KU>B?IUG;cA_IY
^I4]3Y1PMUSc>]82+9L2LM?a_\U#@c.T,BAZB5>Z2A_MYW&P7R:?TENU^]T7^5gI
9:3_^>O@d]dVF37M?Dg0[\?SUJ<)3,ZI#A=WgbH7W\^4BZAXdR#]f1HU8SL6EeF]
S,[ET5HB+ccZJ[^EMKT=6ID(..XH0eVaV^NV5dS>PgG0:0UTcJ+J3FG0;5c.XLd+
G>GBMJWQ6DJ1+^FMU_)HPZHVY_/\-W2KPH7(eM0>O84,<]C.MWb6+9B5U\fO[#e5
_c;\(9,=DQEc>d#HF5S?^Y=/6.=T<f^<daN?1J6-P7O2gf>.SfdN,X34BbF.eKQH
<C^cCL=0R?4[7AfJ:&2]5P3_]dTG6e.308+_H&1R>)bIB(ND&@XA#:N]7\T0:_G(
d@9X>^>2GPCf_>gBg@fONE4VLY\CJd7LZ@a4gK5KEc\D(D==Xe[g]>6/^ed#8S6]
W2JS8#2;@RR1@eX(^IHRPTJ(GR7LV]3)6V1#9D4H+&/g+.H42.]./XV1JQ]<e06\
:&a6aP_c;5UE;7?>&W@78:2IZR3).Qg6S:Gf3K@PZ3DcL)Vg+/\bfZ(EYMGg>G2S
[YbWf,K0A42EGHT+T40:age7@gO5gYMg^]69]O/MCZ/5_21ZN.NVEQ7[_.HG3AW(
PVJa3)>=73]P=T>3caZK51G2L\83]Z<XBHUMTPd<:><J\B;E#d]Gg52B(KRf#WW]
S-+=[/L)V)Me[f,;N@H+XSZJ9TW\GH+HV/4&bIE2_4ITg8N]8F1YfW2M10=5\^J@
-@WbG(IEV>^+D\-<6_aD\5SBZRC/fO0WMM&,0BD?e[>9M^/?@c3gLGXUK(<]RG(\
6+ZXdAJcCeIaRMMD[^7ROGMQK1adMg;M;Rb7PJ]:]IB+AGMF\??E:3F#VY.=^YVF
/X)?I)b,NVaa0YgT&g>/VJ_51YdJ:3PgB?--/73?fGWf5)>6XT=]ae(-1cEI&C<L
JFVd<G4V]=S_B;1;:HD1,@FRbK@e<KIL&9Y/PD11:^YEIYXT]&^E)#c^6If<]#\C
N-VL)g[SeWO^fb:b:<e&HQd)3THe@EWVDOA3>D=SU_SKTLd@ZO0N0V_DU=>ZGHQ7
6J.1&B3_2@SI82\1HU,<JP4-F#Jc2Y+0cC4b4CHUbb]U?G&P0,D^B[:eRd\RG[(a
>4MC9=dbBVC;Ad.C)]+-?MVAd4P?@-,gLG_SS,,2V(GXRRDK\&;-Z8d5N07fQRS=
ec\[K.3)[L/VL<cHT&#9Qbe;KZB2UJ@&aKW73^?+B82)@fe;RQX8@<75U6CI)AOa
HgaQbBM+AJXfIT)EAg77\FI^]J^&Vc@S->gY:f5I7OC^EY+\0[U8HZI8K;b1cI8@
I^PX^9=;@)T3I[d(_d0PXG>a>.YPDJMX7bgAFNK(@/;FHXb9b<7FDN_8Oc>_L7P.
6b^H@e60OgCID5=;K@Bag+WLSLZg\[bL+Zd12@Zg;WP5&SNg?R(SK6bJ8Zc_P>E)
eN],ODN>CU>A-1.4Xg#G\Z+:?eA4g0EG.U:#BV]\DDR0F=P/#4:KF95CX]e;>d^+
Z0TRX\A@1Q_eN)SHdPJ9UP)=A1@?E+CV;ZYX-W7S6EBf;;002GA&g>3(Cb+eK\CS
@&.[7.\Na#MO:0O,&^>S-&/KIAP[fA]IN4I@cBd\?<(25gP3RV#B_KMPb=XJ135.
=0@U?N/(D:3gC(.L,=D86J<db[?dCR4ESd0dR./WLYL/K^BPNZ:D]:8.1V3<V992
R0Pd_L-S:T]Ag7,S2/b#dd8+e](6+83-Re(K;HVPGQ&5e&]GAe&XG3OD#<\?Jeb)
I(RFB_#=ZOR-2Nd>bdW);@J,95NWRR?g0,W)1(5O6RZcZ^9]IS>Rg\4FL8CE,B/#
&=ZN+DB9RT+V-S=+d[(VW5L>7S//BQ2L](L#H;-g,bM2]>.2^AB3]VE>Re#Xg+D>
:JaSDFHf6^-G>U\e-+SDa:B6O-Q9>ZENgFD0(F6)HG0[]&:?a5K]_O70aedPgFH#
\.SPQN-05)RO2?9CLeAd];(U5H3BTe#O8.=>I>f.I4_88Q)0aTCNd0T=.?6QP];L
WGQ@M)R:#Y>K/U0V2\V_NSSeeg^;31f\N/9P0.Kc5C9>V\0\Q;;8(XO=TMZLd8)8
_E,#.RK4:/M?6@QD[V;H#],WK2CR_gF4U7P.D34R?1U2X\Fb+a>44MVObAD8261\
RVGXUVgVC?1UWN+C>-/<PA5N2f?)KU?^DQVA23GT/Ig.\T6)0ZH6G.GN\MTGXY:1
eb:#5+_H[d@&E.c.U[TFdYO3B.;M@URf\M)=2dZR>K=AX9KLRS5@+#CS[a7DT^(X
8/4@3M)ZS^a<b/(X@[3+^23f:gUPBf5KRJ\Pd(_YG\1SVQPK&#2>3;ZHKH&?:0CC
b(=H+(NY]Id,f1ZFMf=S=RdW^205SCTP]Gc1-B7ZNZg,61M\S(KA\U?;F.RH7I?[
N&J:#M1@0]\IVfZ.;aE2+4#126_]:AbWH5RG.SF6-P:cUHBA/CPO=L?=SY^_X1V7
a3-0I9Y4V.ANYVDF0L;-e<@#^Z1a?FW>VE7f6RcFO&PVT066C]H&0G)KM^(,S<3=
.>;>^g_:/<UgIJHCd]0):FdJF1IIbH2X@<WS=RXN(2HE<7CHd?D9R:cA0g<E3f]8
>,f,d=5M-H25<C,eg/aL)SWW@6(4N+aIC=-LX_c=JXdfACR:8568ed66DHTgCP);
UWMN1>70(C_9We<KY\@)K#c8+bVHb>(d-HIW@gK^X2TbFNc<4G-6[L=>8@0=?g#9
8)DN6/2ZJb:M_WW8Ygc]a9E3Y/V.Nb)Z<(?BR//4O,[eLcIc^Wbe/4EP&b_5[eKc
_J>#[cQJCW34&K-.3gE&=QYI?59H,OYX10C77:(b,73a0QdZ2GZ9)DX4I0a_G6?\
8?_J;8Sg0bL9@Q1gO6>N)^<QTTF6Ygf1H8gOJB/D.T2,>JI,41YSLJWYQ+&Ob9X,
f4/^)cU?2&&0B^,7=3+T:@T1LC.L8c8(c&dI<+ET/+8L<_2>L6H(USMYES3.(K4E
Iadg(#I@QOR7(Lf4S8TY&^TY.&H#N9.3M1PTMLG?M:1(g1N#8SV6deOPU)IO=3<&
]L47R<2;M[,21fB1aUX/e1PC+9]MV,EC/c(YA656TNd5-Mf;K3gK^C,=X8X&?0M2
9+QBQJ8V+D9[c4BU_9a1ge4LI_e7>>3)dWabEFgY_=4DSCS8H:-)I]:W?dI3cJ>5
b-e(UJMg<WKb)SE/+@0CGf@PSXJ9dAf.A:R248)_UYf2@NPW\>6bL:^DU_Q6e]=,
]W.&b=NR3N_GHU>Ig,#aAOa[RTfS9e./>aaWZ9e#2_<MAN/-^6a^0-36Ka;\7@Q[
^Q:BFGGWC+&6BJgc)FH(,H\);R-\bc,Z8PV&Y9Da\_E^4KJ-E(8V<>?/6\d4-HXR
_).9G7M8RQM^c2LE>-I,c3Z9-:ZL88E1BA9F\JTJ[=)P#V9EX6A>P_@EBBXQ,48T
e0_-=Q(EU>447<6:ZbY&RWM]43-P]I.>]KI)X&PUP=-<GHDTJJH8]=0V33<4(G4>
C,Z54DE]Ra05SQ<Db-eC\ZQR9\=0b52580>G?B[A#V6:YFC[S,:[FT@92)7U6AK1
\:V=T7ZgDMT@T7e-&(PbUaGY:964-dS?&^-]64fS_:Q0=C>SEBS)^cf[Rc>Y;BCD
<@5gb2<aDQYe[1@GR]Ce8N8\ZC#Y\>TaY\7-c+OA?TVcP947,HQ:&(7V\+=^MRfZ
CJZafaEEg=49J@UWZ@c743(]]#H]F9MCX,C?K<bdA?HOF:#fV]Hb<(R0;debB<<L
dMbMf#DP+P#78<]IYA_?Xb17G=:>2CZa]<TA)cb6Qba[BF?;J>BLcT(X&)ZW04<D
2EKFZ.-72(Y.RB.A2Z8@)K(VA\DFRUQ@N)[F)b^820;52W,X\3aR#ARN+)-?d45g
5J<@58A/E[X+(H-QEF(:U1g>6HI9=<Vb&@4Zc?,e=L[Ug]@3X,ec<8.f@>B]>@(,
_;_]&2EA+e:6WVGag.2J7U+O7f37/I)8Y5HQGDH\Q?5]b1)a;4GPR=68gNCZURDE
P]5]Z<),QB@/_;@29V/b#f>-?IDWSGTGP>GM9Y>D:G(N9N7F^,cfFH/S.WEK\S)^
:PYS(TAK[[]fXc7(@PB?+NNI3>PZO_V0KWC->6MIW[b2VERWB&c@Dg6#9W\fNTV)
Jc[R>@c_D93KC=e[)/=N@M4@EA?^VEdG.bW@b-10271IN/[(N\DAQ+AJY5bM)FgW
T8G-JVd,--.O56QUJdVHeKI-&<-M=K);P/KR](OPT[^\0C2M)GM@(QAe(XHAb^gL
:ff0O(<b)<VRGLS<Te[)NVEO73dRd4.8:VE7.?RK<AIYdN]#B58U:>UZ#D[2+F)c
FL5AC^.a(H4C\25YRb\R)QD@S[T(@5?0_SDcJbN4L/[<^OcI1U826IVN)1L\HL&^
\1f1L^e7EJ0<SA)EfQWc3B8XN4T#OFdedV:7&4Y/_^1)>O?/Y<?)^daTb,L5++[_
@:AM8G-XHcWB?G3K2fVOeWM3L(9e]7]<4V[L@&\#Z[1LCb3.TAHeQKS7(8^]]U4.
.F0/G?IP>g0Ff1<ES^PIWebQVJa/WC&23Z+d2\=\^S/^0@SYK)675<9VL?-YS;[M
H?_81MeC@&^6eV\]dRb#X37:^OQ0b0.(FX_H(42,_+Bd44FWAUZNP78_(B/IXMXP
:^aSQYQU+.R>5.Y70fObg)9KJX0^/OA=gGS0PD]=5cZW[:Og]6^:NbSP_WF=\Y82
X^ZP]Q;&d\X?(BN\2\436QV#?&6;-X8FF?d\B+M?fcdT>>>8d-dSC67\\#YB8(O6
G<^#-9.-?_P5+/H_c\48:?BeeXD3AHfS10NQHQL]VTW3AeA=MUBba=aQK?F<-J7/
A7e13[N5.+1>.#]81FW+@/NT0N3(@>T58K4D?VP/Q\WbWCX\S@I988-2<=QXNgOH
a?;_X@/,&+WSV_Nf)-+>1TP#?Z-.)ZfSF:I:C<TKESPBCU2Fg85G0N0b]4>=KZ42
_1:IQZN&7O+D0\<9Z.);Sd65DN:HQKF4#O-,ZQA()\-0\OVa[#COLPJD57EHP)]\
_<3NG<T_7RS8.++BHGD2YgS87;EG5X0MU:AFgW]QH8e0#VSRH]N7(\[A+9Iff;_4
JQV/Xg4D16ER-JX^@[L])39d(5dH\)J.:bWQF[<)?809+X/X+eMJ\_FagH@S5Cg:
N<5=Y:c&d31gg75(J-BBDU[;/I42<7KR:RB4AadEY^Cad^WET/?+g-#9fTPXDQ:>
P+Vc5dGFU#FNB6Efg+RfB3TffU.QV<0?^6U7?IQ1ZDSWPEQHAcKZY7)1-A75&G>N
dWY3Vb)GfCQ:T/J>#Df4f>9cVN[(f<<S)@d4\(^6G0<He+<P5Pd<L.;RJ@::?TN_
^gJEOE:BAH((b)&O^TF-=^YX2IcW,6d#OAPW7XI@-[VBLS^a9,c9e3ELB+fO_Ab?
G:g@V71)SG/f1PYIJ>c.NZcLY4T/GN[MaWf0(GT;,CNCcGHRJZ1-\&HN^22MCR:O
S=6b=^e/FCbGGD;>G(X-7_<S^Ra5Z]RJD5#KaB0c>PD2]0]F]BK4La]]Kb9K[bLY
38QCa>5]^8J#a3dd=DS\cU/?H05<2?aON=B>O?RNVZ]L5UQgX8R0+GZ.gV;EQU,b
?+/>^&Pf@cLN=.6/.H&F8,6;UA0F8H7J5FTT)9N+6]KG>@88;B]S#_.^1]UfGK,_
.F(gWUeg\UdT.VC>7PZUPWQ\;T9;\YOT:+<+PUBZ/U9J0?-d]P[,;9&I)(FeURAB
gVM-28g4LBE1P.Zdb)]5R=-BL>DHH<H;<P49ge.aJBJ-Ud1W#U(^/T7X+gMHg<cG
A_E(MNag(6X,Kg(;@P^95g\G])BPd\9U8N)+L10Ab,:+W[07feK.<HAXCYL7S=0T
LD@7Ne@c):BCdNc581C-?T&17CV)Bdf&fY2UC1RY25YfaE1KTBG\L^]BKIa=AR2<
0+f1fE<ED+W\MQ0\5<1eTL^DMQ9gd<[NCOLQ7WP?3WQ;4+EJG;=I_d3R,_c7U/LO
@0TVaLZeLM^BWWc:X_PU<TWELab2^,WBPJ,K;\)[[(<CSM;NTAK8BEKK<2-\2g0-
CVc>\WNOET<?T6E>B0\aI)QcfgNKg_cTT7IVMIeH98I^;e?ID;Q<b+Gb#dF5]K4B
<)7V?cPQI69P=c[[30LNI_/:7,CNe1F8SbY8OKF&,eV::\YgWM#bZ-2K9OL,4G>R
cGPNW0e,G.Q-8I)OS_03F_;P(2CW5E+X)IKPWOT&A>:e>_/N)HJCb8]LTY)1.PI7
7W:d7PBP.CKa+.E=G]4IMg=T=19Kg3c,JIUWP+S\+T;+P0</83Q1f\C>P2&(C:<B
HE,La,#V6U8R7IR-Y>/N(QYc5.J6-GB\)TGFB-DT-(N4,+e&+Z527XON),c2Ub>T
?.PQ#N:N4fcH;a18#E&bcHKHcW12.4@PXFcgE#.>IRTAZ[L:cDZ_=E68#VT4USIB
G>48ROJL3EEg;Xe<31(P(#gebM[D7LV4TbTW^,,-a8WaT&6\DgQ:.Q7PN/@CJR<]
,D321#LN8TF.&K.^>EA-F9\LUK<59:N=807b]a6IJR0,JFJD^gaf1#,T:1Q+F37:
eUg)f;H791KGa/(,::N&Z+R:5d_/Q=B=+0?:;gE;?;T<<I\dFJ(e&MAg/>2;TY6-
XC+F.#)7.)2N9;bN4=YP_dN\.)a>8,//.bU[C=bg:LR:AAb6RfR8ZeE]EK05/9,&
JGYF?<HIeGIO;C1(D:\bf(NN+6g31^&?R-\N=Y:gLFg65,Y)QMP6>0[JT0IKCW#b
Ig3YW7C\R@b?&YT@0/0],Q\#FS[(I>(G\<8X04]2eB^PJd/P6F.@HU#R/O5G5MP)
b(6fQ4B>K.=R;XT<BWQY49;JO/@>:Cf6)].gHU3.IfLg7:Gc\fAX72M;DCM\OIHR
NOf7U2c]eF4I1EbM^7L>&=-:N;-(L30(FU:cL)Z/-G,GHK97g=TcLP,BR64@S_E9
B/KITPHX>QZ9+7gM5;IYVadQ2bOLE4KdA>F71R^#b>.Jb/R=RF_A/^ceMZB<<FdW
gC-&6EX<,F?B-PXc<=D\b@;C\V]E+c?QFTDP6DV//B]cAS?AB?cd?Xg[DS[;)(,4
cM^KV?H7<;Z)8[8;,J<9W_/ScaU<V[A;d#S=Je_Bd7O:Y:f>]V\+d1Q8a5dB4HJW
C#^&^@G4GEY?#?dLF=B<O2O0cI<d7HWE&HM/Ec(54@&,:Ra?S868,35MXN[K2=96
7I>4,@BR>>?)()bEHc);8]ML;SMFKc->J6D1<&C60O[eU7HbNbV19/CIGU:ZJDeL
PZ@J4COQ4YW_92-Dd5YY.U,JD.W_b>IJ]13gLEXfLfK).BGNU6J\65+Q.bNEMaQ4
GL6=N^7X3TXU.C]P4.7@#PK^]/fK1J>bb&]OB1b7Bgb4\^,W#G?X:[G]:]23/G)S
0QC_W+<cF_6Y[ZC:/4N<0T[,<3/WW]29bV&6FR/FaMZRU9-YOTb&([a@3#DS_;a3
>YQ66D^Kd@],AB=@XFU,>6Z?GOIeLY&)1NU9L_[bQ/?X;/4B&)6-cA7&f+>&-?<?
6@M.bB6AK?S19FM;]WZMY9H)F@^C?A>FIK7+<[<,Y597;PB(dEeZ7BGUS^W,H-<\
5dN:0a]P]BO[;&@31L/WSPab.RA-CQ)5^EbQLb@+6?L1+^+([:8U0DgUSTJ)gLN5
IC&_FJ>.H1E@I3LN.J.8#cKBDUZa?bLYEU#g/;K+/<FVPEL5,c83?[)HWPfBA)(P
cc^0B+KG>K^J:7.=g4B?\2bODV(.3d@BV1GB8gA6PWbL#1>b8B?=:@BeaN>0LZgN
Vag3Z^)\WGY2/\:bW7[3;N,fCS8U0AXQ]Z71QF.fOO<ABW,AI&0UOSP)I6-a>32c
:=CNDaDG4Ie:X].[7e+KT>Z(@4:M&M:3.W@6KE5(]2Hf6Q__B)e:A:;[<\[&3_=A
0-PHZdKc7G\BHW-c?(E\0:bQ\\9?-K:DT6dC^+L7-X[UQJ:eXTQ@5/7OAWA.FPcB
5QK4SNS3.2N?NE6?HN&BN5+>ZfN,gZMAXfU/>9+APPd5-M=TL;IFMB]bR>_UbAK#
-[c5V,Kf,@=2-:YUae4U2(2+c7TfA2fFSO,CEF)D>)g?U8D<(<=_EZec<)ZRB<U(
HH+@,BM)<DcRZF[HZ4@dCP4&O0QK.1+_+BZEFL28b+)A?HQJ:V0-Pa:Yf__E/c<+
<130MR(XU(,(TgV^ScYcQ.baFUM(g@C0J3[J1D](+c_/Y?)<^T08<4/AE=77eBIX
3]?O&Nb1Y0T\P.3WC\4VeKM(O._],Y:8^gC>1P9dY7gWR\@OSb?DW4=PeQUQ/@=a
dQ)XEXN^0<>\XJYSTW?AM8V8d/P8#d5U5?JZ9@F-J_Z7OP,F7Ee;<)K,E,89>-8I
?S(UDK\DOHSgWef^7QNeLNfHZD3dQW-P4>FJFA28-#A[?]::D&@VZd\1-5-Q2dd-
MUNe>cB1c9P.L](/@=/AF0P^PcDI/LS130S:)[>#;MUY@1M]W30f>aRD1V,[,Xa8
7aPY6#22/a\0/X0Z=\C_B9-90;JfaJ1+3N_3fcPW]#\]X5V_Y[T><cQXeSI[SK3.
9_:.gT3&0bcB@aJZR;TU<gHNE)_ac>TZWS923-ULPA2:S=I5;a6_.=_;UHJ323>[
ARJ[F\@V(W.QbMP<YZ<0?4?(=GP+Ye?]1&U#@Rd]6@&W@Q3;3R5SE@:6:MKA8Y?.
+TB,N9G0UF@0WIB&C<Q9G?Z0:DgC8?@+bgf5[<LTI0_HB(V]0GcbJXR8B;_.fF&8
AE0_f(5[J4HD<W:f:T69+2>^<3;Z-#f;NN7c^#4gd>[?3T,]?(M)+8ISd5BSb5&#
XO,RK62HAB8g.\31Ib<@ccc[UNK>OEZ</E[0QbZ7YfU;R[U[Vc5X?<DJ2G6+B8&F
GY)G0=E:Y:;\>N6@<T(WI(b2Q#M3cBR+eTVU;=<,D+;.>D6AbX/<WQV0<-FZJVB@
OJ&6HB(I@CUAO\[5\7#gUF&[bJSJYd[F8PN@GNB#9JNR-^[5BV?\bT>OQM;<>#>b
HbP-^<9dY]fD>/@8J>:O1-(A?@<0I/?d-;M.RX4M,d,8&]0US?F3?g0_\#<L__(c
@=QFdG.F?XbYcIJ?9e]I7PU_ESXeGDM[b8.KVGNI.(8;,H^_PRSWQMXa2+O\OFTN
[_d&AES:_&-F/W_\8T_8<0D-U.[&1Z7>2>#a>dY6KR3?JK\FedKKS+=3fc@8ZOZ>
4<f-SMZ]C6Y.L[eZ&^J^46Y<T#XZgR\3L,S_0D9X-Zg96S<HX_^HRO],)PQLRL7b
3N)#.Wa)3BL/FU@?-]MNCL]c7+b-T#0Q>a-N?HDWL4VLUKG^K(-Z]&TW@bM3?aL-
&B-/E?1.9?EZD_EGa1,Y8&YBZcIZd^UH;@E9&>\\5Jg:][f-.?ZXSYLL77AZ1+E1
JaQg02FCc#,E=ge6M-81?.eSaJ]?I:@+36+AWM7VV>,_B]Zf_d=(L4P[8D8/NKF0
47\Y8=7NGBaFP5A\A?@Z=_\_f0TU5@1KcJ]C,O@7A#LRgGUBOC5PFIc?S1,3_H=4
];B-O+V2JIATXJe8b4YY\eIVGBgbF(F_HAZ,Yce&cOCb..c<;4bBU_bJH:2T?HXc
??+7(\ecLa;JT)Q19?7D4LY-\@^7]>A34H]N?eS/J@EARgEHEA0a#9.<^,J^4Q(K
I3]Y1LQI)<70S//W/fT+c+(c(L@W&V>=QLMF4)-2bYb0Y]5YPfM,N<6<F:(dJQW5
G]b?YH)2Xb5[AH_BX<K-da)1)?RY,GT<KEUeCIB^\f\Sg3fef9UL_F5F+W[^Yb4;
BB-<2@;H,VYWG+6CfVGgN0Sg1d7&GKGa3f]#O]b?,ROCLD3;AOLTeE/4ZGG^RMVO
5Y7+)>E:=f3<C1/e287a=3cV.4:]1>e&BAe8V[I33>CEA9^4@O(R>_8)g8R[cC@]
-gdFZ5PVc66K_?2#bDXE+9Gg[7[V[#:[^ce=6VTOY2<(8D-Ag(99T&GHNNJ^@\Je
__Ee5dW4FHSRL(MLC?2OKX,Z0fGPcfb1N]\,Lc7,MO32P>eH?JWPNSJ_-]ZX]fWg
:g+GM#,21e?c;B>@I.;[f26a;bP0^0]g0FJ^A,c,2GF1HW+D:-PFH(3&<.cOSfaB
Zce;CGdMA_>ZXWIKF2V)=CMR3W(R;2(M\c:bG-3C2@gGb5a^:D\FVAC>BfRf1]c[
T.D+WODc=@If?df7))W5GAa2D1NS>Q>:6C3<I=-KV+1KOR]/XR>3/6DFag)Cf&@c
TUOH&27g,36>0U,+T^O?JETG[1+I:?[gZ_>-a,Kd=f)YH.Og:PGY5Me2M2W^G/T.
7W1C(XX67EZKACY?U[a)F\H.=ME_3R+SfM75a)XNefIcZI6^Xb32b]VU[:Q49[A7
G#<XU=-+-6)(IT&9FGFZ,[&.E57[H:)/M@9?ED[KcFO9-E^TKUI.SVJQX2^_Z[SJ
Hf]RRL#(-b(ZbIQgG1e:4&C.N/CM8Md4RRaX[K#R,S9;AWG\8+1#,@W/0fCZ9B\[
LacDcY>YSI+2L?(#bZI=CJIZ_J&WU2[<YBDfebc6NC(VHV[W2Cb-O4b:X_JYQ.#E
JT._3:\#P07<+aO14070A=7c<Q3#3OF#/bb)T.=0f@IMd4J?^NaLgS,b,TZ5g=:P
HL0cTM+S9b[C3TEGNPc158\[XaVOabCN(V4(O9IW>C&d#f)7I?RQDW7Gg7UDP^>&
HRTaI#?aPfe67RDN#0>TA<gb;#R0]HQV?)Z2)Q_fB+))f)E5F^CbV043T[4KV)4M
P9QI)69.,&f:\51(@GgHGG(UVe=8,_I(X1F2K@<7J3bH+GY3[6.&5BN->25][\\b
gN3L,RSTB?g=TU1;(7MQ\5J?IgK;^Vfc9LY:C(CL0(->RL(&W:[S,,Y66e6BcecA
>,VZQ/c4G:a=Ce1g\ZK0FXHE@?H^X:I02?WH]fX5d?ALW#D-Y2/YKPG0df9[AL\:
c>T#OJFce@;M&)&P7F8].3S^b?9Z+\cX.ACRJ3#YX#TAK_FaT]XeAXT\^-cB)Na4
:ZXa[ZY6Ra]PJ6V]g5Sa4.bFG51_U1CgBTC^-f\F?116_HH.A?MIPdR0(>KXD9X9
BIZQ/ZE)-XDS\YC&^_g>@f3I^BCAC]d2bgd4VeDD.<0[)=A_7(]N][^48-T>G1]<
]5/QFKSKBf[<4GfC;:T&2b0W;R2J[E/Z7#eBD3I2SSATY1aZbZ?XRT/3#G.D5,[Q
K]8Hd0[bU;fEL)E97WFSZ&OSc?fGLMKXQX4E]MQ,MbN^gFDR=cO:OWJPO/HEY+N=
6A/<RID5a+F<X,?bH#98ODW@?0?@5<IOHBd@(eJQ4Z7EK4;6#3DG5TS3FabLL7,2
bFMg70X42GE0Z(.1^V6AXeGE-1a=S_Ze#WYM3d^Jf9.IPGgeBTWa(,Q]XLAM&b<C
7T8O,L_S/Fgf8CH4-MPM9U.)9G?B.WR\&J3##O3^/_a&DM8#?NO&&?X?)9FO/W+:
XSU>eS)G]LW>TAN#P1H_-N4Pdf[G1]RUIE4gBJ:aE[UV2/WcB>CTgZ)P]COK1JB>
c2]^Bf0NT4?gcQb&LOSCA@:VWLD&N_QfQZEHE5OO@d&aP:4AKN#0?H#@8J^b0&S\
2#C:#EOY-47(1].N9Ma_eF;SGF8GgKE1&cg^U72?cB7@F/S&^]OU6.dR#HbJ6DKT
ZX&M_-X97>I207>R6BYbEfLQcVbd)ad+GY-O,9K[P\SW2.b=+D++3K:(WJW\5_F+
[^9FEMDA<(,5(E]1LA#XGSB3.#4(IPbb7F7+1,DJ;9MHO797JC.H+K_bBPODZW1:
(E3c4S]ZJXC09,_#/D4)N)?JE-#DJ<U+a.adNPg.5g3HVQ[)2/_0dOW4a?;-)P]a
gAMg[(&/H=_PWNA/1W7VLZfUOP+]C+(_43fA29cA=XV3YB/^TX2C:#0_ZZ8Zf1_<
GcP-T.((EX&b2XU)\V7bFL=C32CMA3C4\GUB)6-B1(^E_TPRR3O8?]cIRJOfZ0g.
Z/43Q0-G#+f9[:+3<0<1X/A3Uf&?e>0WB=9cUV21_\LVD[[=,9Rg?]c)-f#d#U;Q
L9IU<Y&68Y@,1(R[BabKGPPYZBE9>AWY&\;U2LGSa]3J.XgK<XS[\Rb8e]/]M7CG
^af6[4SOLVWMY-RT3CE79C2ANMbD5#?H@DaGL+a-BNDF/^]A<0UFZ>DN@gb9BJ/a
62b)Nc15>HP2LA-8Q1)7;]/5\]CbeG:=1BAaXL01IB\I?S,89gR#g;#b83X^#&;c
^Ld^O\Xf(;e(#?A;.,6,OVbcUg1TaV;5M)JRJ(>V>]P/B#W@(YcE.?RO&SZfXB:M
,G\,U)Va^UF?XfeDf8UbOT\=.R.OHCJS<@A#+_N5;;6Z_X7LL(N2,09]SI0OQ-2I
BKKUa\bNH(S^6&QfEabB1)[KYVf/Z^YB]ecMG@R&50@\bLA]Z4OaM<3S)09,695c
L0]a[Y6Hf)B@X2.a-+N:;)19]945\UHe5Z-&0T^T+==X=P)aQBWf)\Q=aU53OW45
<IXfGH1)bX063Ccf3PV5[W\@KJ6EKg77+_R273A:::99e4RP:/DZe1=UKX[9XS;&
ZXU5H11#?_N>E9g1FDbG6R;9B,R=PTc>)9:HUEgdW12#80HX/>GW-..>X)G8^4)+
F8UB#433^QQR&1f\I7BG:FC6LJHADOd2LJ2[?<LNQRZ[5=2J+BNW:L]^ZS2>f_ZW
5\U&OR<1f-&&Z7.L9;/Y9<S]\>eCR15aeX(>HNF;Z\GJag_M)HV08AHdT=/H^^FB
>fc9F,AM18e4T?1K+ZB.dB^Zb6JNAAga=,eKHQYAg@AR1R_,:^LNgI/g23U-QZ3-
19<G\SaMc.<</W;f3?<=25H=d1:AfS[>JV)Ua;21H:J:7XY+OQP[KI3G,QT54U2.
(S_(.QL>FG+JY(@H<:f.g1<0O]J.c4\6N&82QR;XBd+KH8Gb=cB+DIQ],?U,L6:+
Z_2L/PBOgb5AS[^\8#F8^()T=GWP@(_K7De.W@/MBd^2^afSA9)FE03_9=C]a2fa
;fD^XPB0C4J.PC<fV[.EfQP5L>]NP8/4(#T;_PI)4>)7=Yd/6gR,f),;;^Q2WRRU
R.(dQ]@6e2W.U1U;P]ODWf87,6f??AG386Pa^E.AReO:X#@d2TP)-?^KQ8ZT<C58
?gJX7+O1LB#<7RYMSgf@U5(0T2YIX5[H?^\O3A4B>R:H@_Ee>dM]WeJ?;6E4LWHB
9)KO^0O;XZ6ER+7O<J=,c;XBEAL5+V+),cPMX3@?P8=fTTILY5OM[5-b4#A@MWVB
7K?/[+D\F6cR</V[:6^ISd7?UJ+NX[G[C(6&7ffB8H.9.Y^eHD]e]R2-@S3;K9a9
M56N:O@e#:ZUPeDBHVc+,Dd;AC51U,-T.<#>XJZFXGG]^d>J_HIZ3bM@TD6FBT+.
^=^)Y^IS15aDALWdZ=Y0Y[OTV(FO09;6;-U>@^+F7S[ZG-T=DVe0E7)?;eQZcFg7
PSNND==.>5T48J<0HOF,@.=JF[b=]a;7=]CG.]3NdQ34VS03D7/B_0?9D=6UD]4b
TX<AT_H5M1JR-g[b(8D2JPZ6[;-IMKATEBB]TO+#;X74RK<W2?9XF]f#F5RL(4db
DT[Dc\:+,Qe+OWTPe#bMM-CB+;-<]CgX/\?Lg2T.;RMQK1E97D(=+<Q#JTUOM/#7
ZQLT#=/G^3L1A[S>5[8+0a9\67,S(NaCM0BbNT>)&:VDC,V02N5BE[=Ub+d2[CE5
f&0K-f2f=\eSac;]RN/cB)1J2ZG3:<-gU0H7<:8S[PVd@8dfWI4Y,P;>PDV[;?^6
+5>JLO^0(A5,KPYDD<<.0W\]@4X#S_VLc_1K.#-]M3M&15-Z83dZDWD2:VJS1QO=
d;ZS#/0JQ+=d,3ceKZ<X?C&=4+eQ4D/YF.6YZ;W.>).1WC3&SY52V@=)>f#Sb2H2
dY_;K6]=gc1L?Z>3cY;.(WKO)UA^PKg[CC2XY75dI_f:feT?eNDJ<:1@L#>?>F+6
>H,VJPKG54c?5N2N?ZOI\E-./XW8]]g4)_MeEde,>0LV+Q1TWYNUGFJLC+](GK[[
_0V;?e-TKL.P@(0.#?IX@DF9K[.=A@K/Pa@EAIfdV#2dJ:TL9^bT\L<,1F]<7Gc.
770d1Hd=28],,.L-d@UYVI;BX3bE(gZ^RNA3628a)Z^83)]M]0,C,cZF0L:D8)@Y
+d66[_^OHE89If=^(OZW5<\?b0[f8A[_bUg_L+T<1EG8(&T<5WI&=LBKYQOH231O
=+UHg0ETH(DK2Gc=]QE6SE.cA1JQ4QNUB^Z2bP?UZb9ca#/_W=GN;eOVacD4:>eJ
#ODH)Z5QKE)G?HW(\Ic><efA5+_f6@:A-/ROQSOO8TL3/:AN1#f.T)O694eW6G3]
]HCC^[&agd/SNW>3,\9INLB1^E]:FWQ@0-&Y/d]H:c/aJIgGZC/[68C_((NGB6bZ
_@&;e[;SW&^)OLX20IJ.\f]b3;\g?9<_Q2E@Ug1=g1+4W3GQ\EUMYM7J=8VZW>_)
A:[:e.@VV6][LYX1H./HceVLd0e5_RWg0\7JfBUgG8MAbdFScTMJQEECcdd+LR+E
-Oc#XAYaaOWb@KgYc>9Z_GKB>E_:9I51LJc-<#=N.Vg#0P:002DeQ#.3&PF50#C6
J)07G&C>4a9OXOYZY^+[AC?0,bD0Q@4;_5V]B+U>5:2g[:aTTF[3IQbf3ZbfYRdb
(K#MDZ)[DRb/M=H08=Rb[Q57+AVP0,>HKbTbUZ>Z<IMG_LH:/\U\B?-M>5QN]a\4
EI.=5aRF23&SD,Jb00Qg6f?a4bOXG;)6JG(3dZK_J9QUGG.=Ce,S3YdQ,^SJIaW6
;(U5H;PR8GIRJgB]0:5<baP5e_ZgJB1)WaKEI96]9g7-H?=ACT1fRP/8YTPS^QfN
e-;QeRAQ6&J(I1+72GX=-J-7I;5NG50<ZF6e26W6eWc@bOK5Cg^DbK>)U)U-13S-
)W286I28M??R+\MF2N>5c90de6Y3,6Tg]Y1TMN0fd>d:=cc,bQFdW8HVX)g_>6=)
XMS43e^,@+ZfD,Jcg/-MT#cTN/DSQKOgUV2J7LX,2E[(,Uf2SL]BN6NTA^87?_/4
c<=TL?/^N/b+(DQR^<&&a)TXPcPZD^7.cf8W[+/&(=cVfef5QS#Q&_F]R;.PT<A2
#4d(bEA6^,5K#+8c1^>D3gAL[aZ&Q10RgSSL(4e-5Y:MAGJM;9eJBg,:GQ4)@Bg^
fCXJMTRMP^7_9ZF7SSS<[TCg>D_,VP^^CI?L1+AKcLU4WDLV5KWR@9WA0fO6?1[V
<ANbg^@<G#VL(SFEL_#]FV8@<VF-#eP<Y&aR#Y>ReL4_F(C[.)F9cW4GY&J?.XW^
\Z.L.b1>F1dc;09;Fe-GL>UAL1<=;E6F-<J0e?LL.P5/<@UK7E13^G##GQG=#(PS
d0f]ICSJA^=\eRSQE.ZaQ^4QNdBcPV(_SaM8S64K^]SX,fK]4C3U/bC@F+>LeJf)
JVUHIP><B4M)>8H40TgFb1]-7YDX@<,LFWV1g-20@GX@1f0gJYEB)RFU((+f1f3<
:Sb;QgM3=9JfN((F2&0:&Q?7b2_b+fQ=K^6LX;.C)4+#9U?>H@+,1,76@)OeNU9^
5Y=3^56W_0^>]ScJ6D03Q:O5,,)X8bG>@b]K;;=&bcYUT>@;2Y<b7//B+:cfe#+O
K6O[TU4\W&5.X\ZX89Xb3.O9O&P9CE3GbQZ&UD[Yg79:T&\aF-:eP=3B(M8<2dS)
aR#ZPS]7+DcG_WM,T@RES-4C)^d6VFIXDg0TVMf3+Ed/F?<MMNECVZUM7_IB,0B?
EL<2[<N7&OXXTPHB3K32E7?=g?bCdeEf(#\d-@#I9EaBQ#eOGCd]G?W)2ITQJg@0
OW(LO7<T5LgI@aI+1_/06+:NX.-M&_4>eUJ?2XU0f,@_(36::)L6E(fE@QAeg[IQ
T;5NQ@A,WIDf:KNF4[>Y82-8cW=;]\d-JZD)b[R+-fa51#fNG4@3(]KIT)(_e#V\
bLSZR-]#?e^d82=CLN8,D7cGQ,_BPQ/2(DC73b&LVK>C4>3cO6-0^f\6=YJ;HC</
./cNeS]BHWZ73c76eEC2\?;(OVbG;>Z_-DKM+d=BS:(ZA#_+3[.&EYfA)cK@?PU&
CV5?SPe#W\,34_<T=edQ::X]BB.Zaa4&Z3_#ZNdR8,F^-E#G;&1Q#0UR\Kd(F[QY
M@WN)[7@^g+96<X,9VP)D>SLDbB61L70R354CN#7OYS.3cC68?QO^E5\:R=.?g[\
a^,?b./bLK)ZaSdA;8IDQ-cbceeL_\BX>=EO[8.,Tb)#[7W.U5<>0:P0f5S_2cG(
VE/G1ZU39R+9_S/1,]Y<PXe].(\.HQZ.&+BQ/BVdQaYL,3I)49VgCRYaD-DM,8+6
(._OH-:D=#:1[V&.:,-R,]./Q<S_&O.DN>T,0fE(+Be+;-fe#_/\eH]/:[1.aHbX
CG^:KMDf(TEAIK<D;LR?\>5abc^Eg9VaZ0aUVgXA9@2(E])6@HE8\B8MPH)B+US]
IM,TCG5E;-^BH:,RZ6b?Z<JRP(-]?QQ>X1Y0W#1_]<3\5#f6Rg;/DS>aM[M0a;)[
e.>65#^3c=>V-UPV_aRMKF?1\e\MENK0/GO)XB(4ZM]H\T<(83UO==OEUI+aCUTU
Bda#J^58I(_HR&K6)V+]<[7Cc=b1E+O))9,@6eFfCec7F+#_gC5#^2c=Bc]8G1SI
X54XGI6I\1)EI:JW/PIg5YWbQJ7ZT,Ve;S/&2;gLb@a^06JYR7O]QA<d>-R890>+
RdRUe7#SWLJE]^([REO;K8(9SAT_1G72bL/bU^6L<1&H+D8_0;,UXAJ2,MaA@32^
VE;NFP)db&R#SY;DZH[1G7-N>Ec-Q8gNBD@[A>,<Z)YBYXe8=K/(VK59VUdPd9J)
039VT-F7PCDe8(W/6e&:L>RW7Xc](S&@HOA+,+JWJONKQ=?g,GNSAJLJ8F<]5bfB
5T.4S.M23^6:Nc#T:Ne(gG;KESZbEX2dIA@X7&3S4C5f;T@M1>aGC26S07-I[#?^
=9d:We(_DXeYMf5>]:G8D;FWUI7#C\d9-8?(U_gcfLC=TPJUFUBZYEOXF0ge(bIF
QIJBO]6TW>F++JX3M5bENOGd)8>0^=QTDT?g-ZKKd#[>Xe)AQIX;O05B-YYcC@K/
XX>J\f;E.]=Y3f7QDB+gRIg4P(JcAe0T[8EZ)_ba>LO-^Kb/Z1G@P\CO4gaO]&5)
X5ZRJ+TT0+J/fPXBEc3[>C+bP.<63(.QLZ?dTAXM4I5U,(.0)4LcW6)@)XW>=\<]
M2gbUcF]L7\8CW+dA2H-C<]SW<V@7<eN4UdcMDR/eIb.NO2,MAZBUfPAQJbWYTRP
]Q,BSaL4g@_9/7CeY(T9=eQ+8@-gTVa27VSKRT)L[+=TMgVS?2fQcT.b:E;dR>UI
-_ZbR?-6dR#M4&BXJ,C+X5PA0<f@97Zef\+^f_F5aQ><@-7.eSE.bM1^CcYU2dC;
Y&4S(4I,0H;O8aFFVJV8d:OA:a2KVbS9NG:eBG0(b3+8II6;3Te5US:g:W@BPKJ5
XZ)UA/=C2J7;c4D^e6W6ND?(2a.e_WOD[=^=9AY5O9_[WB91.T4TE9^IOVZXdA?/
U:HDCF&4LbWL1NPcA-JeQa+^WUZE,8AXP3\ZXU6CEA94aJe8]4[BOM^28TX5UI8>
@-6<1;5AY67=&=R=[RGQ4)ABKJZ9IZ<P/G/WS8Oec?GfLWURRKXCSHTd&#E@:aL;
^7K73WJ\b&<:QKT3d:b\KO]^@cDTfHE4,C@Mf[g7UED,W\)CD:F[#_T5P/8>V1[N
c>(H.R+54.U>,a9E7?_MeBg(?@8BQ+#,)/O8H&-G6bD6^.DT#+(X5Bg88K-A<ED2
-PbB&N:6AA2_O3N5J_SO795W_E]+_<0F+A5(dP(c6PT)/dTI@[F(DA#?QYK.BI&J
<6M_LGWBYGMWc3M_Bf4EL.XC0,O:e.>VGV:cV-@RHO^D4HWPF_Xd1>VYbTE/4a5\
DF/Y-PPOC+D1(5:=Z;P@X592+^K3U@@QC?VU3&YcBBf^+?\<afA0VY<?U\H\XDIL
KTI(K,2.F075?TLW.A-_K1d@UeKB(2SF,307FHCM;-5c/[@9eUB9U7S4E.9=\;[b
1<8Y>Z#A9CbVeSdP77dcYSTN_5A@,9[2&gY/F]WTX4W5K&e\<+:WT3L?MeS-2JSW
O1B858O]@P.(#;9BF04EPM7I/0A#O]_M+dJZDHR[=J8c=,:P1?(a\\-g2S2N:fV\
_U][>_BO9UP6SNfYH?)]TGFU3Y=@SO,MQCFY15K+N((-L/=Yfg2UCOM2W+1SPQL5
Qa;fZCGR2bIOVV[>QUR]C_5\2+Q#,4\aFa/INb&6))=0@VH\L-L@LBLOA0RYEAZI
:fQdX]V30=YA31@c\Nd/aKfCe@_9L=1=]De#IaXg8CZf-1SUHPGU.[Z(-132NQR6
<@d@Oa8f;823Q[c0He9_;-_=(XG\HJ+:[01C.,Qd=P-QTBYJc4B:<c5/7#<0C-g#
[?2b7BXO3/Q1^TV3FT-G_+P[N]?7,+[MJ5S#LcXWW#ZY>VKE1SYZ/TD-P(,NKC73
T1d-CI9)C^0S^W5V12QQaHDKLK9..gZSP8;KIR:H+5:1NK2UE(J#CS[^Q[BM=YAF
=BKJP)6-TIA4EJ2L:OOb141R-H<??fM1GS3X)DYQfd8Z2F,HMZC=9,W:HWa+:MHK
:P&QSfN]PH>5LN^MX:R/(7KI4@LX7=I)CTb&Y7MR>RFMcZ.J--1B9V#8O3<16BS1
)QID#Z--9ZS@<8HIZgcN]NBF,L9)RD?,_?CNL)5fba9MNY2CGVT&YUJ@_OXb\3&D
4P?U_M0=6L24(0BP=OTKe;#>M.cH;g=e/Fb]]a)1b37#e&g=V)Ea^RHBcJ&?0SL\
FKKXU:NB>F@].>QF8BRV>92X2[NcPeT1MCaBdCRYM1;fI@7,bd.SX&,F_#F:TN(/
F8K3K_9OQECe091+\XFB+;a)J+#JcOQb<3<(N+CC0ZETCBL_<87Pc,c0fgDV7(W7
gKX]<,N+-.SR76^NK8[9,[Z0<^>8QN-2.>T96H([.bYac\f^Bg>>EMMR=&IfYeKD
GI]#g=6EQ9JR@Y@HZSWb[[F6/P_YTDSUWe/+?NgL__)#_23\,E^GS-:JN:OC#B57
a:HPGIQ:,Ac;8+A+5GN#J7\b\ZC-eWFcG\?<:K.^4N;V>R5_,#EYSC2;[Y^T4.\J
ODg.cEUKbUIBSId504UHgSH/Z]^_]>3]88FI]&1DG#\6<)_VEeEIX:VWHGGE:>#2
UB,JH/H\)+aRe025X\OC;Z^KS[.?&KB_+VJWH:4\GB.B+8)+F&&XORZ0ZKOP0-[^
T>48RdZCc18M_e3V;.2e.+9(74Y>T0f/X\AAGC5+@c8=-GL:C.T;a(bAZMg+S4@1
)fM))YDIC.]VQc143_E_9/.&7C4=&:>4IBMNTPG+L&0FL-S:dcZadN0gc=g\W0cR
>W1=R-X7O9OKXUDHXKX9=O.EK+?[GOKZHgI,(,#[94IO2OV,gNN(?@IcUX[X:=9+
JR7,Y&VRK?W>EYB?fY&]<9J0[:HW8__\FWgb0>.b:DLUE_b#0[I]<RVc?85O=Ec4
Ie2?E11;PY71V1K]TJNHO_N@PW17):.YE2gbI<J<M)3RROE89Yd_7<62?SO@WAV?
IQ7LWW(TEZ7T&CGMc)07_[IA[3]O:K((Me>Y8+X)>cT:X,SDBH1K>]YF1@6=:,JU
1T<^HfWP-PQ?6+bBMCT:,RWQ_bQ(:d^L-U5bQT\9ePK];Tc/D)?6\NdS62R<70Z&
>6FeKU<XfW[;)862,C414-de)=3T#YGag37MD9JV6[f>N:_\5gZ5=SgI_0E9=Y4Z
[)-=S&dEVMeHUJ5(YRK)Z_<U038-(B8]NJ^:7Q0g?TMETZ>-H2I90SKf@946CZE9
@+[3FKJ3S60MV\)#,+.4W4/9IG-;8S9dX)_5\:af?:(#9feS_gT-OYc9&c:M(IO[
U8?T8b\?]eW,7c[2JX4-+-B(O;->DWM#4?c6=+b/@44fR,M(5&a[I98SEVf/I([,
aN70_3c&V=CI^g;cg(gFFTeL\F).DTQLL7N1QKP<E&Fe.^Wd2FM0TX,86W&9WZ>#
/AQX=[=\cYS;g8X,M855\C-#@]ffI>CT9<&L(R,PIN]H-(92<WW>(=V#;OIU&@X6
#DE/Z2).@<98PZ+6(IdaK]g6)(<09N[fZTP86dEGe=9G(CA:LcULEe<1d[:ISKD#
30faAA]N0DY4cG??N#JHg,#9GH&EO3?8G#1567;8A8&82^VAfMXQO0H[-aA#-(#L
Z12]7)S>;JM:MJTNW@_6c.VI/^ZV]A##P5[Yc=f,-TEK1KW3&1546bYc9:=4Na-<
a;ESKN>PdZ?g3MbQWZA5M>E>F3M<8+b-I)HP\ED(a.FW8=7<X(K\[5XU8Ag3]3R2
K0^G@4S54,_aBS/V#dfg_Ef-OC&;RJW+>S03ZTfSMS@F_K3:8[?VD1GJf(-?E;2[
-/TES(U\)@#L/=>XP-?:N+KXUc>YS:RC])ZDRCgC5?TgEG=T8=.#<V9N03==TOZe
Z]8^2gN<bdAXQ_>-H1B61Z\V@J8S>^9N\9O;)&YI]N_+6[BU>_#F(QC@QV8C-bW8
:=3F]3afe0R[;aZEY7;3XR5M?Wa\&Rcb#_gD?ZdOXHWR7F^TJ]WW3eK)\4O-XK>9
Ye7bG]Oe)SB=2[6T;fA723ObEXZ6K1PgFNaD?B?]C-I+DSQ.?gMK6W+Rc=E0(;O?
?OSAeb@O0L#a&;C3\eLUL3YA/OCBB2A(,[LC@=<Z83\+9Ea?\^eUE8dDZ[95H3?g
H:,\2\+X9T_5BU?B84\#Z</&V[ZNZ0fgVZ[)ZM9LcGW0AE]>:>]#OOO4+NM3;b/Z
\,3@==]M3cAIgXY3@cPHaH+dg]LWEQ:XZN(I6NYgLMR]L;4<YdV:,&Hcd()?VQHK
3WI9g)>C++#&eP7,X_J#3:Kc1dMgaL<@T]B3I^C6SLd\FgYBc/JRMR^:2QUZKc-R
aT+IOE0#QdP#N=L71.cNTD\V70G&]V;8aK.IWb(I@QDON>AMR+Q19(?.KRAb2.?,
6RKFBdJ>7S#.eTeCF=?SMa6:gPF\9:<;e(4FaS3XYJF>O3]X=<4SVRF:Pb/VSVI:
[.]RR^,bB@,d\CV8Z(N,\=+O_7J]Q3e<GU3g7JKUQfQ;P+PGBNANQ\UNeXMCU\@:
g:XO0VdZ?.V)7#a(-&-.K0/9Z\9D3<=((^PTPJ)0]]TZgdgKV5gO+1aTM&aD9=LI
<G60[E[-6.F^@^<<JBef9:84Re7]aa6W-G.FS,\f?XcfV;M;Q9C;^O#P&@e^A18/
XM1&;/#TCKSN?Hc4f8SXKf=#EH^-J/&CaGed40RTSZ9M_:XXH+43GE1KDH,.TRX>
3IbT#W/W(RKff:0R^J-]MLO:I65.US#QS\7X)OQXcSW:_?LSg7]Fc79ag[+^>QU4
H.-3N;0EZa/N53gF,P[#]HWL0[=aXO8<e_B90JN&G]E[9SD#cLF_^>P^:EJAQA#U
CB>FY<UNG7]^d;+K60cgfVP[@SEC6:NQL3<bRLGE+=(8_W3+EM]8+[U.&+)Sf/<d
b67M7P;3Yf\d<0d5a,2=@,4&:0[^PQQU9<79\29047-REUfZ4[NXEb\[6U=JbcWJ
=DV27T6T^<5DRSDO3Ae2UI:L07S^Kd(XF5X4>@LF:?3+cL35/4d2HQWF&3@X>/Yd
-18B4U&=/9IRLNY:[HG1JaDTVXJDT:>=VT:F.MH)GdcGG\(<Z?;043C:30Xd(0cE
<Rg7K(0M-De)(HH1eQGJXT\E?f2=&91D[5V>XH(-(+M#M_gJg6&Z7NUDHKAGVBg-
g&R4BNdV>/V[@&1?b</]I:1SS?PW(.V+PXcc&[X0QV2.FR])8]XJLCA&-<U_#<4J
S3A.P[gUg(.d@]F6RJU-[?QeeQMa)Bf,eb?_c=76^UNM>^2O_M=;F3G6I;5^+R4c
EUJ:PB656B<OP2Cf3QTB@J]g&f6C&I7fWJ@IeG=0=#5^9FFQ9\&&fXZ[bDe^TYaL
_CP)AA][TgRQZ0B0Fa2B9+L&M_PF1I5,8)Cb3Q):0bK,T/9=\U0>0,dS;.77BgS5
:EXBcKa@GLI0MfWN1,H)W3I/R[[:OW0J@:I+>N(..L4g][FXcRb;Z9FS^,^).ca9
-dJ)VI;L:##eR&)fbb2aKRYQK)FR:.<L<-?bQO)1[gA2N[bcg,F_CVK=dJMEGOMJ
94TRDN-(V]<+<[)V,VBc7#(DMJ==+S0eH@3,/O?Xf_@/9@NS0Nf(XR7WF.KN0XSZ
<R<^e>&f4D@-\1;<N58A#65+8J:0eWc1ZY>)8<98NGIbC<A,US../@9b>/6R^\eJ
f^K/O41VOgAc\XADT4HUgSJSHGY,J:FI,VU#.VZT4Y[6;8;5&SIKI,I:LDJ.K41@
66BQL6M5T)<O,TM#MV,2cNS^L.1(5)gRVK.PG1FP0JQLF;]5^fa)YfPJ:16914B6
7Z[DW)3#^<^GAHBGKN:_WdE/Y1PX=?EV/=O^aJ1O#FW2H4;A/718BbDU(bBV<;9L
6E9bBYVddLP-[)@H:Z8,M6FBS4_<O&-aCZ38LO/F,MJTgQI(@DU2@(YUH#J_KEZ:
D>R/5g;5J3&Q/Y65,Q=We_2MfFIISOOgZ9aM,[>bd.IFB,XI[4:A7V/^LW0J?26A
JA)&UBN_WI5a\QRT0,+T1E/(6R:.(NcH0Y87B+(X1^?RHL3N_?.NC<Q5_^B+2-1Z
H2#:E97f:7K[:6KYPQ,8Q9-W+0K,OI\EOWe4K448:S=Y3^d[M.DF(\G9HAaR#,=Z
E;-GQ10M[X+TP+XH--b5@/X(GIJ&#;b3C#2N;fBZ6O,BOG-dYC2XC(eXNKZ.g6Ab
;9EbIJ4@^6R@F9RSJf9@cGD#N#&X)+R>([^6<M0=S)e79.\U+>E>T?)Q==Y^@S3M
>]@PW68N(8(1W9MX?]/F3b;FHA10?+H5(QK7[3a++K(E(XI&JZJ\<J)>,A4/N(L]
_,b</(5^80&691LBfSgJebR7b5E0R1Rb@/WB,02FJ>HYX&AMFN\fQQ=B6K;A1J=R
2CS8O>8<[b@UY@DI)T__;(72<#RIe?D9a9UPS^BDNP3D1>G0/e:[;RNHNNaE9U6C
0/&dH-9gaRB8ZU.c:fNF8)K@-6XUSU<T^D,2ANe1c/8,Q;f_1CGJ:.?\[N&ZX<SI
dA6YHWcPX:CUBMP0OL.((6Tb6F]-<OW2SQ-:Q#8@f(2;Q#/9_S>Z9K>PUf,#_GVD
)F)?_UA+EgbQ2L?g4@IG7;f:=N=Mc=M-[B=2NWLcde@1#ZLaGaIN9H930Xg,>(ND
dUK0D8ND-C-+-eE[FPMNY<&HF<_-W2]8^;TK)H?7OBYgINMMSEF-f>Y(9X/F>RD9
\KWW]J5GK9)=T=DD;Pf<gHC:+B_)UAHRV3de=B8O[;e@4>/]O,@LOU97Q<BYU,-S
gf^@UEES-3f0CU\aTVXBT=QP2G8dQBG/)DO]VC#J6bP@1-1I=SG^g8T+fPXf^^5d
LFb(XCK)T9+QY6Va24=(JZa&ZHAdRgT1+#O#8^M5R<@>6:+L?cDc7fbC;Q7UH5QT
KfN#7JdK3g,Kd;B;)K1C\b3LTY47FAMF9S3Qg5gf<3:P[/K<2&LP(MX+acbIR:T[
HT;OTB14?O#3]2B2B\,3Pa9E<95PK03W:UXAL9^E^bDA+JGR-a9;_a+)[SOK2Z9B
_<U6G-:@X9YOD-Q53>[AERJA6a(9XQQCW9U=Fe+;eCB82e&_3\3PEf?70;QfcF&R
c:R8G,.)(@S<9[9(Q?<A=_6B7VCa7R8;4g+E&FKVb0))<XNMHM)#0Ec9?+0cC/g=
^/#4e]^S\K#FPDIE:<aLcFDS>GXgS7Z^5O&Z_DPEEQ-L3HU:=\&J63-U7@&XKac4
CN_XJO\@^Q-#B3cVg-T5[WZ0+/eXba:0L,R^PEH@VdBX7)GD^:W[B-=F6B#5Uc0?
.FdMAQ1)cdXb5=[JKM2.U#c\0aE7b8Q(U6=GU[D3M?NX<#g.]F]7Zf@O?58fJTX\
CM0ZN\0\T3,OgU5BAW+EP-B=[d)#S1>14=^@OS=U/8.WT/V<^?9C,T[)[9(Ue7A.
L)-=B@91\5-3M]gCfI?I_JYX@L==1RU_^\2XA)8WA,CI_;;gWW1+>H^/EaT,=BY^
=:.eS,c,<^BH+OfL=K+bd(_Yb;dE.W<^:3]3cTbS&ASRR0&3P3Aa-g6[>T8]b>UF
e5Ue@J.X2&(,Sa.C3,B\J]DJ[[IX&+->cZ3a;8B#=[gHgQIdc>DaYN08C>3UcIFP
4LC<CE#5Y&dZW(]GNX9X8YNK8UKLeG#G=?(,99cJL(c/\U;8b:S2])JN)>(6bMT9
c6KX0SAP\/P[KA45,V5BC)]I)+)C7T./5;(cUX?K55\]7(:?R=8#/[F;M?b/.5fe
?WDS@>\-QWP[RgY7fXBcg6#bb2W<JWMR1\@P_O[FMM:=P_-d>F6QB7&O(_R1ATGK
:AS#>J5GFb=)GR3UB=62GF,@JA/XEI@,MSMS=#_=468]5<g2R2g7E?PM55CJ0:Y)
DaIQ&W@16g74Na1BJ<[)@]V==7_M>/GG1_.;NdK5XSZZ[HI&_=^Fge;U<F^A@K_6
>2bL&)M;dKA-cK(?PAF<;?SOH<_gB,BC<;b#]]c&4bFN+5\T?J^ZR.a:[NPU;@8Y
B@>Z&Ua;==@OMZ?M@C,#MXg2-H(fD0PX#3/?b.RZ9A7E[Rg75G8;WT>@XT3ED7Ac
8RO^R8L07+NS]=PT8bE;b[ff7Qa9K+V\gB.L@F0aU9aDVA>>3#CfeNJTSCBgLdgR
^dYN\E&VM@L+Q;SO<)U@&@a5SN66/2L7fdZ\0V\<+=JDOcK@9f9Qg43deKRY72J#
bgg5&YT3JJ4RRAO.QS5PPA)3OZCAQa_Q@D,15;VADI_6)025O-NICZ=f,b.G\BI:
669B]@I[\?\a\JI2OW&:0aCEaK#c)LV4RD1,bFf>5fcFX-\^68/G@N\.Q]^C^_D#
BB1G;QX<RdP@ZS[]1C-?fHU\[H/YL1XXec)Ud&1+P#\e_4Yg64APSKBOEJ^4f<Za
cfC]&W81f2PX>\WU-]d#508+E=Z8F1<D6ag\B/bZ=XZ+_-(,557f?NQMg86+_e6W
\53P;I[,C;B+_+<-7CY?2]<NM(5CC2=^HY-\Jc6YDB:Y;d2KEPND].Dc[VX\37@2
-&,64@S]LgZ[+[-7+]78T4\FZfATQ1B?MG>4<5&E2Le:b[[RKKddVb,XL0TM7KDM
-.NS>RS3L7696R@0a@+7gH>Z.O>.XNE43f+YH.HQEQ;-@aB941VS3,3e)&b?_5C;
.FB35>KO#K1;W;>:RXVIT0@aG3HW#0+S_KSFBS/bHHT@/<:7RPE60[4&XPcL8UBG
\WQ&-&]GBVIO^N#cf+0==;B]W/(3</\;TQ6,L8#D>R>KJ\ZI7K237(C8G?c_bMRJ
QfDadd[?;WCU;Z4J^aa@gc7([[:5?TJL8WeNO5)2fIUQ+?[R.9ZaT_RIM>/228I5
_LF6fDQJ;VaQGBR=LgJ1M(<_#)K>&P>JC0(D)&]3)fY.JNV.c0D54f&,<b,:6f8H
bdg]=P>G^?F]]4VQ76[T?^P>/]:b]7-a_gC=K\A@9C3J:]cT_)Uf.F^8G<b-b#-D
KZW>(&8[GA:a0JBI+;>3;QI#5A?#_[Z<K-d@HP]_4<5FV-f\efged9>IHbUFI/gH
KecI<K<EcEF6d#c512aAM7BMAcf-C&2]&d5I>+SUC?=[IT)#09(6?))Z1SM9&RGI
N5fKgWe#L<Q]RB?&-=H?ELS1-I6N8@0_d75FD)_b4ZMf4c#IcgKgB,;a^#Od>.5H
H=0\A0S0E/V3a67;THP3K)\EC,#Ag,/X;_TO2NJYSSIW80X<_C,R\?WgYB.1LYeQ
Vg./5#24eOV]Zeb+R-)#LE7FLGcW4CR@U5-H9X9NCP:3e\f.d64C99B4E0)[cQR[
OS)U@;0<gXE[F)6?g8,eb;Ya<;DOgR&F7DVR:=b^TIaLL731a]27QA\87BX^#6R[
PT>E\8ePR]aHA>7gH(I3H<Gb-3WH:BV/>(T9,69AJ]aaZ-ZB?Sc\@e/C89Tg+>Q;
ga:]P_9G:ZCfBAI-/2[>6BW-RPU1_>2Z.]AJ)NCSWU.;VF5aDW7FMSdf8?;e]1_T
?6+T[MOI:37TX0H]?D_Z/)#9,NY]G3YR9JKOG69NfLe0;+g=fe-Q8?:E#Lg;6L5]
d-.#T?)CTb^-XI:41++[XL]gg@>+G@38>>B90U4_JG;WHX>DXK_L.d._FXCT[DOe
93dYH5A/XD9SeXe;P9@RITA/??Gc&M/bB06;cU1bBbMQbULgMCST7OFH.RT2Z(+c
\^OaSX^_Bd97?C6e>7TXXHb:P6H7HY4T;ZB.<O2\@^aBa:.f/35+Ib6^#e[RQ--:
E(F<.Oa,PLgSgNa0BQ:8Ie1bYMPL-8/MXNN5NP.]V.C:3EDgELEZ8?I()H]_(L-K
DELcce<I&M<SJEA;1agNg,JF-ZUbC56J)E02=cLT^(R+.;Sd0A((PP_=eW&@LL_Q
aB]ARgbP7P_()T?_F>\D8>+M)01^6HH.MgeZ;QMJWPHDbO+[\.:9;BFDKNQD(8U3
/27DM<bCUWM,bO1H^(N[PGdO5g&Le9=E_&7J(d9V?]<aF.X>d3a-W>H6\gf^3#P5
;?7aab3SWS#5_?dRN[[V(RX;K>7IRa=K4Y<fA]745,5H7bDNSDQ4SQ[g:48:FSDZ
J)G+9D]Y))+R;PEFTbZ3JJWR2<^A+&J&eRdO_76=IfO7>Kf&B1^L6c(K6RHE;?7Y
QY&3)gL=&?.,3739I]ID4G>1J\GE-J00A1Z=OZ80^,N4_GeRZS2eX(#1Ja26c2E5
a(ecRM,:96779(XUY9OCL[+b4.4M[c+cBA15\U\L=Z8;]IO#8bDVTLNJ.dKQ#bD)
HW7eKMQKYP@U,XZ&90?9AEQ0gW^>PX@\J+3O-ZCT-X4,]Sc#@B&[W(gd52B[7/JP
PMd+#IJ3)[S:\2KEeM1[-B6IX@ELG>N?FZ2D8?:Z[:-cDRR-,HYNSO.4Tb)[@G^g
;D;[[0#.6=Q4a@>EeWB\=-a-@MMWQ,-MT653MNf]0FIcA+&_.O0,]35Cb,.NGdX^
K/LV[IN&8_4^8X@NVN,JK)UUff6VN_YEE-S>FcfOY+RL_KMeJD.Bf]:HCaBJ.g?M
UW600Af;E=E=4)+>cL;\+?R;]P-/D[1P6MNO\T2R=)1(6KC_WFNY1FWRAfBX#DH(
HM((6[6T#GG4..=TV5f>d[Q>FK\ZCa26ZIfA2OAWc\]fKJRa>FKDO(MM9Bd=Q6]/
1.Ec0fT#&ec)4&3E1#6D+J-:4S+7;/+.#<BT,>\:c2cFSYg^c2c[;2\_Rdc(R)_,
?S-U.VL_(&Ud?Q6\+cfUb=g@3E?<IJT:7/T)2TbBe4>f;3(Z>E8KC+4AeJ>+&K&R
<F/6U/4-U,0I4_NBO1.?Ya2Wd[1N7G#V]3B@]VMXc/P14H;&&LX0<.1Y>gH03fW)
DHP8&(]7(O:+dUY:@:;bJJfYT&GT;I,dOQKe5WBg/(M]Q&#7;,+?1]R86>#O#5\0
gX4^4;6YO[Hg0F0^5e\5c2fU3?F<;<fTBd#YQIYGXQ,,^^f/A^\]Pe247M<QSNE?
2]^6O38GQZ;6&Y#,PcEIX\E<?;eM?X;Z?2IacZTNZ&.dS5QU]c45EGU:(9#;3AW@
BB@;:L?]b&=Vg&(I<:TfYBS5,e[\_IK=V,;b>F17#/AI0#8H0H=Y<]/3/QO:[7J9
#6+.0.L7_TT8-YR7JZR[?HQ?W14aE9LfOCM/A,Q/G(:WQ4>BXQ-6Y/65TE#JU3@_
^PXTa2\4CVRPAF@#4^[]1M(+9\)bg([OFZ+6-]=MG#/3E^@=:#Xc.NC@RAP)^bP,
YA<ec\M^([6;AMQ>SOEQ70/bd]+Zf&N#U0J1\1D-NS70718a<J7^FZ&,RB64HI99
WOOBI(1ab^dG<7gMgNVY@6/01:L#=_&081RA9cH1SX==\;3QOU&C?(T60JeV7,YR
C#YPOM2cLD:c3(JFYAL/f<b#ZR9Xb)<BAT7MZ_1Bg]S:C2K=<TUWDM5Kdf<NJOd2
JT.&eN(W6E+<J>552dZ)8U)4I^,fT,AA+/.Ee/0)#5^?=^G1[BOD:(GN2-Q3K<A6
C6NdX^V3B??,EA3PDK_&;,g8VZM8L+=&J\@Qf\H2I<OG62X<ePaEOeg8(Q^+ZXc\
a/XJR;X(4?b)I6Y.A^:g:fU:M8()ZW[.SRY5PO(SG//Td2Fe<BXa/AW)[MYfEbG#
C.ee7=FWY)L9O^0GbED##aEKHMb7C6f]dFVFDIBB\MQ@/3W24),T(Z=D??Z68;c(
S@#)e6I^,Dg7ILIcH79#?]SN3a:H;FV:D&+1ONQ>BB]Ma-OC,-MR,YNO7ASD)4OI
L)d<eS^6GVIRW9:U,DL/SJQ]#4+7E6-\25<6SWg9>U6O\?e1Fb0QJ1Wb&AT1:cAR
-@G3eZ:1A<T@K/6^^W6I;d6ASS=7a.^U?R&:aX^BL]A-]<+X2DDgfPI3P1;#3#P1
G321B\+2f89&AaB+VaC>:4(2aPR(O(^cI7,=J:3#Za-U2[L-G@A5OCTSU.#b((&c
?2aKZ,&2?CTSe778ecPS4G2+C0GgX0LW(S#d\KV;<gD8@>#\DHJ3cMWMd64,BQW^
Ha#e4\_7GLH#NRCaW#ADR1T3_5YNU+F8,PdQGNMW,P)<f8+79)eeGC6&VLWC6_aQ
F2RF=.(5?MUfG<b,Q93\25Q23Wd9?2>:_CdbYJ:DN=c?<EPDTAD,2I_,X;AgSEd8
QXYLE>Y25Wae;[[I,OA.<aG#;<=)G(I)<XZ70_5E&MK0)cY8IZNK9,gUA^NC8M-D
>9(KGa+CVQ8F92@a]ZOMX2Z\(La?S8P3F#WX8ggc>@1.a^427\c<(_#,b3+G7=1Z
PV,AB_ETN^Bg+/6_FC<FDY6XP.NZ&CY.+=FDN&KeK4Hf=,-FE2,[2LH],^c)_0N^
-\_@,.GYM6>-)PLVb>MW6X0a_8^QXG.HcK>J^=[,#-eB(ETf<]<e(=,F@6Y@f_VX
?DfG1]CI+1(\B.#9@6#;X^0f\Y+Lf3eU;;ZdfDS,C#0;HYYH=9Z5PH.=7:B[=Gd)
a[4g2J;NH9+P&]7>S19);FC(7.;4/7&K+Lg:IL#-#+6>OR&STSRR8a7@VFAZ2E;5
D63X(MLG.2a6=[;NZR-(X4NT9X&8NX/8ZS1&#]9X)QgLa]^#,eAI2S&.a[Le#e(G
+1gbW)_XdTWFR1-(AOU3B55V121B3/OY2RS--[V:TW)U^;Z0R1+^HaL[Q4JZM==H
O@GV#CXDaEGM[A<=f(g:66c?Ve)a^D8gWO#\d1_0(?<BI-d.TA.eH<X#7?_MbQVQ
^^&,(ZJP1H=ZFB++OMN9X[?PS?P&Y[bF31NX<g_&58J_SV1[1#\WR@B9[X/#ZbMA
)BVZ<T<,I<5]??ZG2F3LRAfL.[dMe^O.efQF1EM?D?5+edT=_&-ZRV/I2d#JK)7U
\Y))-gN[[,+Y?9e3_+3^[MR4XOJcBH5b159)^-6N7LZN4XBa=?])X[9FNeNT]>-M
Z50Vec&(@-2YR#]V=AO,I>)P&f7E@_X;Ze[ReP9g3aLMPFgIbd8O^S4C+XWS@UQU
5G<Yd9.\gGbI>X/4Zg1Ke\GLI[d88PPZQc;],gI_X@W5(Y^R<\3WK2dH]8^S]1c8
^b.;[(SXJaKEbH>&:/K3+]Vf&C@DH5(Y0_XSA/<T<9-QG?(Q[+0Fc#Pd[D.&g\;_
T+^&X^TQ+><=;P?,FR[Y3Wbd>1^7aH2/18<BacC1IdeT)G2#_gY#-DR0CcHY+Xe)
(?TKP3(<X&TUL^NSSN[V]Mg4[]4=7;.IE3dd3L(VJK?-4\;W_[?b5#TJ51QFePP?
WCQ^7C];\(5bCFIe.-,KE]fgO\c:?JX6>718^4e4[ZQ6a3^ROWKf3d1cf[L[NK#7
D^VUHeFCSPX4+KW]cF3ZX?e:f5b9P7#_15HX@55GNL61L1:@#;]5d,QFB5P)LaC\
BMELPOCM<[/_P;>Mg+=-6,HQUM789&b(=NYBV6S6>_OF53>YW]YA=Id)5eLVC._[
E>#AW@ZE>/-A[g\[f:3<O9_a6bWD+X\JDUHb)&8HU9ab7+H,e^(3AJgXKOB@U?D&
d183VDVXA3GV<4dZ_7B+g4NK/.eY73^D4W#\296?5E^g&:>BSCf)MLE6X.C6\2A3
P]YJ<DgT4RNa__RO+dBaDagDV1XU04?BaEbZ9I#VT6RX;KR:TP;Q?dECP2W(Nc[6
@5O_1.HIF2G8(-Y:d#99P+B6G2cY;J]RWZ^;IS]].IAIgZX(.47Y/27W@HGFN1]_
5@349Ba^5-[(@ZKfGabdQF8AKB4C&L&#@0.UFg>-P9c)[(QfG4Qa[L:S&)6H2gQI
I01FP@9[@7)S&2MMfGdZ\fP-R\IMQI/\O4:#G(C@8H2-Ab&9PfYXDgNN8.>,Ac@_
0E1\^6MYY/:b_IE_9d3GFOL-AZYYVCB_V;2;_\Z?\[/BE(+^#6(g9MCMZ8)?]E<E
WXaD\ba)bU4#2[\1O0L^FRGB1fRI1gWdZfG(+8Y+R>f#S67_A#Y0<Z+edG_cDb#O
>\DaN1.SES>I-,J.7+=@RU<ZPBS@/VDX,XQJ<5KO+\ODJ-?7G_P;-g;GC@/]^;?<
XdW/LLHK6P)Z9f2N/NLR9.eXSFTbV48W1[6,D9?Sf#c[DD(:+;PaPH?GJO_SNM]0
03#20e3/6EQ\RG)##5ISX^.#&.#LU?70H-P2\gDT.NHJU#0[ZU)/+_(?]9g(DZ7-
NQ0/4G92U[4O]GW#<bfXfDR])OQD@3SU3WCMeBO0YW<a,f@W]gEX?H@_<P/dT]ZJ
+S_4F/SG?AB/MB;K2;;LgG8f[]].+Q0R7:C;Pda;)X-(,P&NfE\eF\1JTK14f:9<
#>QFJ0(X4.G_T2&S9=;a]-9L]C[44,:XN1cNGD;Q0c/3+<LO?VP0GRF=&eReO(Me
;7Ya?P-\U]FPPd>UbcJc]CJaVOL70I8\g@&+3FCDaD?,)5Y8A(W3;AVR2]g=ROR?
[F;.Q[GQQRXW<EYIMB-MN#,B(6:c3d(\EW0L;74->Z5A6[[ZfXC]EaDUE(F8.&Ig
^=0@RDcON)a.4:]X<HODeTR7L1BN@]e7]Y\(:45WaVabA4LeDD=T7NGA/NU-^E_,
?,?E;.L^@Y=08_dV0Rd1&eR5a_fUg>I/aDBG#Hb8&^BU^9_8b8NcK4g+bP8gJ2@a
GJ1^[\e_3C[,L:e@7IWVf/)_(D.-YPO&7F6/GK_WWIL[Ya.:6@>AGd]?K7_Ca[a.
?<##CNa5Q>DgYPIMJV)\8Z>7]GBH(\53XL=NRHYWLceG&VWI7P+g261=Z>UbPc(d
_XVJ[J(\[8#6/:Jf8f7]LZ_=M],,.0:SZ9N]P<I4ZI1X&W.<)W:#>7.(?68-f^d6
7(cX,>A4Da@R00Wa.T?JK<A.cbQT71L+QX,E18AY2;#>+4^Q4X5.O6NgYW6T.O:L
S>_I0S#eAE))CQ=+W/<.@E3GEA)E&M_QMG;Y,W+]3]NGe--.Cf,gN;2&_0?8^M7(
YUQ;JNc5W&@.L/V+(_T>N[?T>P#?T[JE]3)f];E/N2MCg>0M3BX^&6Qb=bH2YQ\P
S@:1)c=[\aX-(:Y/;[2cP(>I1RQBRL+gU)(fN).XL56LW0=Z,aL#9g#1B;fZ>UCe
1PA:6C,H1IeBR8+1K9LDcA3OHH[T2^,F+)0c;5g_][GCE]_V:WWWbT8[DQT4X3EU
N(bAW+,9;?#I/FP(SKS+Wc;7<P_[?)dD]JP],EV.OYJH;6XFZG9,GFc@f_OdS4/1
JS;JLUW(.K_f+5I[=G?-c@E=:Vd0c2d:EC+M.8&ecUFS(/:=41MM6+B(bZ8^W--6
X7Y+KdE<IF207D34JAS584PN65NX0EOZ?;8(J\\W0f#KX#?875[0JY+UBe@)P1GD
e8cc1eYA9cYP3@b8c>(6fe[/>;eQga5Nbdf<6G#F,VKCdN(9=;=gKMN7)VG1J5O^
^P,NeX(53TT3,V7(_GZS4I816/]9;H9BVc75JNd#M.fV+(DF0GHIIF>4@GZRB_2E
8U\^^4fLVXbTP6MCU6JeVO@g(/)-J<QEU8g:P>f5_[b<LC21Rc^=VXFZ0LK,EJ5Y
7+MPQe&>e>M)dFCL&2+4A[:_)fDS5QR9D[3M7IMI]=B-JQKQV,4g@L3Q>cRQ;R0L
URXI<7>^KOL[U)YTVbK;LFI:1gad#V1_EFB&XPPfc0L0H)6Y:8PESN-8BP\D#[IF
MaMZ7UK2;JHZN)b_fe+MA_VO@^?cL?.X[+GgZ2JW.L,+g=32VE^2&ZT<((#3cW26
JA39>\LWUX+cN_-b_J[1.e0=_g6=6/XJ\aUf[e)GWG]b-XGIU&,@^f)@Dd8.4__?
P]Gg1UWP\MK2IWe,QJM5>L=L,gedA(RJ.#4TE2ZHVWdadGLcC1KVV],;C)dS:F_c
a_Y)J2QB]a)5BGQT5I/9LZ]-7NLK4E(G.#K&]LQI,@-ZQ@EBTb3\,)JJAVa9gG&-
Ja9caTD;Pg@<N2-I@0cG1R70H#:4=MQW5]<8739P\OK74A&V6cEEgXC]E>-c-c8_
<gVg?XB@=_X@(57B[JA7ZIB;(BcJSBV.aE96G-TcQefD69_Z5I<7)9JP:8JE_X+W
E;?9@+LNJ;+PVV-Aga?G;K>[/]d<<,(4;JJ)9B;(eMS&F@L;#=\Q3^:[.0Z7(H3e
A1bLW)fI.3Ca>0D-(^gCGgEBg(aZ5]Xc=Uc&MYd)6-OC<=SFgE0=@2gVL/>baB1S
Q[AMS99PA+Q1F&LL:A.fK7ZS1S268.@<Z7,L>I)fQ-a)0f\R[<T0KHgNgLN)\;.P
T:,51JfgaA>g\DGFJ35E?3[4gJZcJ.9-a4\f^;ZG)&eEGe@_TQd(EaKUN9A0b9WT
IO@e<@&;9>4=<UD02YNV4Q+IXMa(eQ/UV1#aNfeaV\;aR9@<(+EP(BU_D0<gU&f9
?g+\]OJH,0F,]GW\E9GF^CB_(WYO[^RYbQCXa8HJBR<]deAQU;,eDLT?<#?.>#7F
F5[EQ-6I-XH8d]5E<C(AKVQe)gX]c:aDT/6NE5Y)da3L=6Z4fIDT+=&-.@c(-0(S
G#=b.OY+VDF5TGc)7GBKLKX1:RgW?eM;U-=+DY\D[+]N#O,B?f5Kb,_g/R+Z)EGL
de)6OE0V.bQdDK3eQN3bD^-R+L84?&T<0QKKH\OX@Z7+AK9XY3UR0EBM8-\ed:d]
SX(U#-J1XdPXb2cDd<W8_6M&De8FM0Q^MedYU,&ZR#.60<b]Sf8+GEIaY(]A43_Q
P0?3LdC6T@7SV3YJ;9P]CN/3DfL^/B(4V1PT[dAFO4>]Y[aFT4W;f&e?P_7,6O1]
)PT4ZG@WJ320#\90c&Ye041fA0F3,PXX_UE\AfMc9G#a;#]FcW5GG6-]&bUHR)^U
5RD#ZI(KA<7O,3,>E4X_TSZ_F^HIAP[9ELTLa8[ZbMHDS/QdefI#ZB-7QJ9T7MH?
@RXfDdX@AB[V(,FZ1U=FMMBV+YB+&:H,>VE1,L2^3Q=/K;5>A<eT)AW\8AO9WHLM
(;7;Q0cJA_K)Gd^=_([#f7a[bYW_#:\Y;NOCdPTBH\BN&X70:<X@1.KVFMLdQ=eE
3._#J@Y?5=?)f8c<aE/^cHXRO81M?cR\<5H8EF(E_[2Q@_&)SZa&:[?_QRT+G9LB
_FOUPaM\2NT)@2f37NHb_#H.BO^I,=K_U&b-9c-F[R8\;,W9Qf\@T<9)JW>[Kf5J
C-#EOTYASGD51UU#XVRNYHKa,8#gHZ1UU.<#TT<+3?\IKRJ)E5VF4Z.INPgVVXWZ
UXJ.eUfRINaNH7NF4,]3?C9P1:S>5gW<.G4VC[>?<O\ddU,0APO<YMJ)D(#S9I^9
P0.K:U:YI^K_H][GWY27C9XY?^Y:9K?&ab16M-RM/S#NYZ+6\.N,3KN])[?gA3<#
AAT86Y_J[5H-V]M;3_aY^W[^(2G7+(a/0f+[.1Q.^)cH.HUQ+VW)@FD[@(Z/N/Me
T6G/\cD[e0UK3;I80ECfE3]>bG>^\PLY3]NN6\#E)AK(b=Dg\]g4R+#L5Cg[?@/2
b<LMaH-FLFFALTAaKcObVRB>eN@RL\Z63G]>:9IZW3Z.;V[3-@442M3/#^/=K3d1
R\]/E<E3C+c:DYJEA7_e]NeJT/gd+\B^_?F+87BM\VMH13HGX86@f],1VHY2]2(U
;;Q7@:H@G-VQ@8#4U=CB7QCVRR>AW5Q>U1(]QOKb00V@[_(f&<.MgO&0a&M2Rgg3
P]SESS9)EJ]]-W7aB=2d^O.FdD+4fB0bW)_=f1/1][L<J^Bf,-X14P_9^ABXd0PZ
\I/#G;?):C0-D4R?a?:/WJQM?[,QA^FC82Ce&Md\-JF<@BNQ:2W9<4Yc9+Z=^?R6
^ZG./-LG@;Y;eTa@,JSW(D4CA#Z)HGJ_M)NOKgQPCBc2PY+)L6_;,K1K3N?NXLZC
NI0(NHSJgQPf=^TTaH:CFVQG]J5M4Q_3Y;M,O>;]KBeNI(_F<?ZF;(dT7f]XD92E
X#N/D#(XTbWNV/P&VZK;fL9&dM+72]7e?@\ICg]aRaB@H13RY#92a@US#8,.fIV4
6KIZAc<e8gI0ad?G(XW)19.f01W<@e)aT>a#ZR-e5(^X)X/J)R<1e3R&Cb/IP@-A
TMPK9:29c@OJ^5>8D95S:>,VOTF3MW(QdUS=,,,:V]SfI(EYJNDe9Y41FZA?7WFb
=Y>Qdc6?AN-3d1Sc9\b^P:F84JQH7IccN8G5\+0\).QTT:DJ^JZ#@T6\ZLS_UXc-
SP\=^fc8G:#DU966<ffMcD;d_[IPTW_L51;M:J]K]=38QZU[bd:fbPc#Y6CL9aT@
ODb+=c\J:6a[UF<NQ(d-+&TOaT:)Z)4W#\Z[5PI>]fM/YP(.W-JGNS;OJ>R9cYe3
Y>5gX4HOP1680.@<FN&gDYagcC+Jb5#JA8d-f3,QFY>9Me=^K?K0TT4@?4RaX?=3
DV<60;MH]10U9VdBY+.7>X&&G_H:D8JSU)NgTP1\B?&)ZUg<J:]]XI2P4@\gT?_G
L33aC7[ZE9-NPIZ@T<CX;B(BY5_^.+LbabQB4\fF473@BTC&-J9#T]Wc0.B\28B7
]E\6Q2JP:S65GQ_dRIgV.>9.8IX-PA)9-C/9N>MM8Q#GOc;Y6:g7RfHBgNdEU>IR
@0@3V\T9fcUAS5&B_G_WG+&fCaD6g_)R<T@^X]+>ZS>_8eI0?S@DYV7R[13]8g+B
-Cb;fbX^X;2g&+]TDP\:MI^Q5O?4X6X:\X,3P<YE.cWO#\g=Q+@/[QbO>^9J19@L
SR[478L0)KBb>_CP97?I>[=e7<8VQ</:D)4I.JQ,UI[P)AdA?fX01J<PF^ZF\\ZR
V@PbXf.EgbW=7_D:Z54R2ga-8H>dMIU1-)GG.a<_cIEe&GY=YCH>FFA;&>LQZ6@0
[bP=W(5[+ILMN:-VSTT(@Y/UUTPZ3gI7WPQ/X<.US@LKZ1O9?d[d;g4\<TW4G6]f
FRDfEC^\IZ-]^5WX_P/9>=2W]3;C\+MRb+IcC7=Z&A=Q?9N7?/FY/5BKIJf2D[TY
e(&6^DE?M?4,/JccRR9-d0PV.K1=6E9#2C?J:4NeR?_\24AQ2+bebgfRbfA7;Q3O
KB+X=gG2aHGC+d^d25WWfLREUE^T<&B:8/TeIg\g16fP1L>=f):IC2QaY1JJ,LgO
<D[1OQg^X4#X\HQPHM.#0Ib0VPWW,^;JXSaY6?^?2I)(/]J6SEQSGP0\E]K_MAeU
P8cC-5bgNbT=1T++SbI?>\TL7;-OTY3c)ga<Z^#<3]DeaF&feHdYP_F=4DOQa+IG
[F5,69O<L#\F878I._MGVID,JAQ41+WV[D2R[MV6Y#\,7[#H[W)3Eb7KgXVdX]Nf
,C3b.Yeb;:(;#5<,70a2:7LIe^7YHLa(:&W)R]FN2E3TVYDG)9<C,CggR>6OI]YC
<^95ROa=H<)[I[3GM2B1\YE?7Z#?Ae)ccCA;(BFAT<NaVRW?R3B0,a2&7XV.3c6D
VJJQUc/;6-@Df/QS6.0]:,(&g\=>SNDL[Z@4EM/=/X)ASKX-NZ8GJE8Fb?=:/MO_
ZX23L>+C=20.gdZ:@I_+C3bJ_ZWZ[#5AM0PXI.UC5,-HffNcGPTU+K3^TF0<Z:G9
>PY#CYB[(.aV(e25fD=ZNfXbH#+98dMMT(-VTCZT8&R84PeDJ9=Sb[+5IS(L1)@>
-ZD9Te@EWYC?:(-:(_P;L?#J@9)]?0LET#\<Fe:d>4AJ-8RYPSDGL]fNO<KSKB?6
bR4#,?K]d.Lfa0#E#L8eR==<,=)28G.S7&;:5_)/MgVAT44J\Z&f4.1)Qd,#\XOB
(b:K\P_5Z>0OC-Z8\N2R?M2HCd3B(\-0Q.b7(=bScfgFbY.7LA^?^RM5P89G^+aY
<-cee&X_TaA_ea,#UF0?Y&_0A6-X\#fQ1(4KF@38Gd)f?IK;YC0),H))Gd+W>d\Y
;X>A^MIafd25=XHG8L-A]OC/,8]\\UQSY@,<DA1:&+2BLXa6DI(e@Y_YI,ANT31J
</LAN=SAF<T.XAQQc@U_\?QCQ;(=b(T\<E1&LRfWVKH?.NVL=#VTB2N9;^cJTS)&
6##4)&(&>K8YP@bL1;5PO:S3dUc]]T(A/Q](#M24&U4;cG64B#IQ(WEB6N;g0@XB
JPB7g:GdC1&gO31)PeHabfJN9>B8TQ#9L#e2B9?&PT.P7):&Jc&RB,-I;eR;DP[,
[M2a+C)XJMgW_KL2Y=IaOZKICc5G3+<8VSF:;Bc:>P&^gY0be5FXX\)WZDc\:)c&
T-^J>eHGe[ee<=fO)FB7J:S/WC45O;E([)]LaB#A]OgDA9d)5R87KSeY8#D9e#Tg
Vc,\:g(#@]aL4+a\#DH#O:P4?d7AOcCfTNUM1-dbZ@Qd12,B9@(-/VR130D^A2IW
RI9;ASEA?UC6R\^PD5DR??W(1=aZa+IHLQTA^acQO.I+U?M+[QLY@,54aK9O@+B/
EW;1=Eb9S2T9QC7=4=KI4A6gCQ4VZ)()=_K^A<d630-]f_/F9U996AUB^4[=e\)^
K<eH&g\F/dA-6Be6dQaPA@9BNb<>bE-1_AbGI<ZaJ8R/SIb=Gd6\.AH)K4/QW2F8
[34U;\_-)7^&S_Me(&+P;?PbJ=g01<:\802_[8ee9b9[WMf>-fIgeVcg8.F\B<PD
1#Ebg1g38.Kf?VZNBIJ//EQH33Je9EMB.&6He>@24c?=SM/e#LAa?K>GN<B^UO^2
?gWZ8S34gHSQg9.GR/APL5f]@?-b]?aB?AC;TWAT3_U/GJ^5UXTce^B:Sfb[d^1@
Q/5Q.6X[f&XMB0EFY)0D[HVQ+Qg76e5&-dc^-Had6K.W9=Ta6Lb]edWX>A3(NC>J
FO\F@eIT&._28:-X/V-AdY]6#]P+FGaUc)S9NF(:eV<Z_F0#?RS+<AOaON#4MdL_
9=J#4K+\+0aCJ6Be:KF/:Vg#C@;6E9,-(V3#2;P]9^&[[;,g_a<4RMaO;&8KM:KK
e2fL-.0;78[K75GCOf:01c:G8LT^Yd[[M1]M[+[INc&&aafaSP1d-E8T2G#L6Q>5
;gBM&6RA._N+-[PQR&16V8Y-)P^LNF_DeHV-Fg..WU=I0P_c9?&]4K2A@;/RNN]\
;N]LOG54\Y640<cf_I1D3G.;:-2BC5;;TTBOYNHA<7,Ja\.g7gO\2b,P<G2RAgP;
MS^P03P3aK8D,[1\@Rb5b7f/DZ+=0#F@[PPI>>8<.ef[JRG^=)ES6f32U3-1A&E:
U+IL)DEM^Z#T2S^cG9R-S5g]5]=deU2SE]ZGBPP<F#b)B+EHH4E)-a2I:gI^ZeWU
EU>P.OWc[_.ef,APaM9JVWY)c#b)B9:;=g8ENT6VK@(D4)/7E#c@V92M..G&-8bL
Yf[NE:7&dEE#cbdd(dF=WGbe^+^SYH@_0e;RAd\E2RGFA(1\S<GE8F:e4fP&g]4M
A?Z4[XdJ\YMTY;:CKSF]T/GcR[Sg:_0BR(UV0^U3)\D&KU=?S@9PKPaG/4[1RX7H
SR=NF2^9/gHc9\5/K#7@PQ(PR0C2EHTcZB8Q\50.dMN5VIS)63d,4BfgPf0QHB48
26_)HcXaf5LcZT4V5NSA;UGE<T-+I0&dcOBb=:cX[dQ#6Lff,aO8DCZ5aa&b=Q+X
,(7#-VVLXJ@<JB[D=E>I9\Z;DdQY#[)12HVf5073D/PA(F#/5_SZK??R;JCVAZcQ
065AR4/3=AGGKf+Z)b_M3g>^V0/O-bM9-2Q9B;g/V@MEP6eFc[0:(O/+LH]JB;TL
:K#NQ?[42^Q8cPeVJ1E:76?^DZ,ggCbZ@Q?VO,&R?9Dcf5PNWb1UK,[4\#N1=88c
d4.bV4]HU/S7eURK?.-V>ePb3UQGaCCA<B=6e[<RQFa9a]b8CU<L-Q4(=IW8>PI;
C-Uc-Z@YQ<Nab9&WB[<KF,dUL.A/O93dI/Hc8[M,9?E<5A>.f)W0W-;AAY8<aDMd
<#KXRH4)PfZ:<P73OVTN;<Y9Tb,G1a39JG2a@;K@HWQ-(DafWbcUHGB0KA&&;Be0
#;67_99_;T3+65bNW7M>]bS9ga\(;F^P&A;M/QMX.22X_=KPLK:=>L<>c8=Vd(>e
/==,+_FO,KWHYZ(a<U1Y]f.T<@L3DX7?\KB6b2Fa[e=S@G;D(&78NdC5fT8QL3LQ
8[2[WQ;N?B0-38Q.F[&G1SG0HNZ.1<K(BO<PGIT?GFA9CPF/QWHJDONeKIe:Ne4T
]?IJUT4b^>GR5DIU;-B.b8HAN@4O9-(O6#TMcUYI3(7:cG9E:]7K#Y6W-FTDJN)L
c?W3g0DYe=^>LO&EZN0Y=eLNf:A2NA-H6O.cY\E?S7fYH(+P?P_[7eX[.66B?QG8
8F83CQD:a&O=KUUH\GTP.]A0=Fcf8W<R[P<dZX#M[=W4TL?E]^@T6C13TZ2(=O([
c@P,QIPD/G=.[81;VDT<I@YS1f\Y4-=54d]c=&=IMP0e+7KRNA&,F?78Q.S0W>\V
NH_[0(.LN?gc+CRW:XA^]C)R3_b[bd]P;;H(D=EWV2+3#,QfAaH[G=/?6:,S?bWW
Va&(RSV08Ibd_<=>O#KK#=QI&D,2?WDFO_-K6]7b0VV?8H@Vf@Z44K#\cD9A(]IW
_9([6e@>&eZ/g\]&f1NEDXX+O24S]?F_-Ob365eL(F)R@\7487cD,7Y;WV\VE9K+
SE\,(;8@CC+]2]<.DZO;+U2JD:gGMJC>>O&&<9V#UD/Ib]O8eWcD^14\;6c[b8KZ
JMG+#(b.gTBB4d8[MQM]-)C72_UUH>+^GafZWI3FX@WNa#@@gV9Oa_B=2f9P,D]e
BE,OVS/E_:c8/3603[dV(c?JR-,4#P:<+8C#VKTU/68R#EPXYB=0?2K7:0K_?dUA
T;dgC;;16.ISG:.X6fIB?]e.-2(4JM2Q+c;(NX<F>X-#O(61)=1Q\[H6f)[-bQH,
76TU+YET)9-cGC)UL0Ye7C)V2GXWLR2eG,O]g0RU-0]X7(X)fKd-_]II9B)3?;3_
..E@G(2T+FSPZcED\6J.;fc2IcH\#0f#PI?5(Fe?_2PZIF>6(H:_bG.22^ZAH--2
N5O@F,A@M,.HWIg/=:a2HKb#4gXO[S#HE-b+>;+7fAC[D\8YQOK(=AX+1^N>ZY\Z
;29;;U&XLQPKcA(:b9^=+G4OB[FG8L)Ld<RLQPELL7+=[E83^+R]@3L]4AN<EN)+
CMZOXV5E^=gYOD([ggefPI,O3?,6?=]PJ^RF+:T@;=D@d]c_,d@0WR4)9MK5g6_#
b0M1&e[-/a.-If:4;&X)A^_4O]L@5\Q0N=1QU@c<P&E<bdc]\9[,:J_FW,IFa3VD
5c5A0Y(,>F75@N?#=QDHU,^C?SX@(YDMQ9I(<H>60A#@;^..,JMO(&9CdCGDS@UA
/b^]LS-a^-^Hg7=;^&g=7Y#:M:g:PJV)X;>9cEGYFSER\77.1BS@D4JW7N:Y6OeB
T+Q/6bSEFOFHOe+/BQ;g96-1[V44WX6L\>=9UBYPI+L>^I0?7=PDb.;fG8D\LSQ_
J<?c4HNe<L_0X&J.a.#\>10FKPADf&7DXReW&gEH91eZ\fPS0S]bYUI)(#VU_<<Q
0?>8-+9,K)(E-\>_cMfVORF)UcVHO(8(C=>PLHNT#6E[>YO8D:/NB?O[_UUJ<af#
R#RfYS5#69FD1.BD&3WXK)X/.J+_Y]-e.0YbRKTTabDRM>8QR9M/\:SLGbMS8LSG
FO(DQMS36VV1ca(?A0c1eA&/QJ71Q7Nb)Ra-]L)EVO_0>4CE/CO7K0f:(:D;=P5F
\,02)SQ-0S=J=@V<Z9HS@D3b(bN[QP&:V(J,)1@Z4=&VB1QLP[d37g,WaU/I3AB?
1fbf4U0-aI>W(JMA5;L7f,OaX)K,fX86C\R<0D,P0BbPMK>ZKFW5-.EA<b^9FfIe
PUQIbBBdL7I7(_AGc9B@a0PA3<;7=@Scb^Uc8U8,aZ-K;P@:e6[HL3/TDU<TUGD(
^2@XcT(R;,RLG&<9Fc[W(48DR2aZ)cJ>/<OI=54=EF&KA$
`endprotected
endmodule

